VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapper_sha1
  CLASS BLOCK ;
  FOREIGN wrapper_sha1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 1000.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 996.000 85.470 1000.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 4.120 1000.000 4.720 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 264.560 1000.000 265.160 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 291.080 1000.000 291.680 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 316.920 1000.000 317.520 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 342.760 1000.000 343.360 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 369.280 1000.000 369.880 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 395.120 1000.000 395.720 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 420.960 1000.000 421.560 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 447.480 1000.000 448.080 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 473.320 1000.000 473.920 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 499.840 1000.000 500.440 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 29.960 1000.000 30.560 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 525.680 1000.000 526.280 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 551.520 1000.000 552.120 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 578.040 1000.000 578.640 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 603.880 1000.000 604.480 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 629.720 1000.000 630.320 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 656.240 1000.000 656.840 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 682.080 1000.000 682.680 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 708.600 1000.000 709.200 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 734.440 1000.000 735.040 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 760.280 1000.000 760.880 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 55.800 1000.000 56.400 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 786.800 1000.000 787.400 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 812.640 1000.000 813.240 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 838.480 1000.000 839.080 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 865.000 1000.000 865.600 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 890.840 1000.000 891.440 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 917.360 1000.000 917.960 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 943.200 1000.000 943.800 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 969.040 1000.000 969.640 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 82.320 1000.000 82.920 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 108.160 1000.000 108.760 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 134.000 1000.000 134.600 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 160.520 1000.000 161.120 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 186.360 1000.000 186.960 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 212.200 1000.000 212.800 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 238.720 1000.000 239.320 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 21.120 1000.000 21.720 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 282.240 1000.000 282.840 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 308.080 1000.000 308.680 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 334.600 1000.000 335.200 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 360.440 1000.000 361.040 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 386.280 1000.000 386.880 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 412.800 1000.000 413.400 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 438.640 1000.000 439.240 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 464.480 1000.000 465.080 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 491.000 1000.000 491.600 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 516.840 1000.000 517.440 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 46.960 1000.000 47.560 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 543.360 1000.000 543.960 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 569.200 1000.000 569.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 595.040 1000.000 595.640 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 621.560 1000.000 622.160 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 647.400 1000.000 648.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 673.240 1000.000 673.840 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 699.760 1000.000 700.360 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 725.600 1000.000 726.200 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 752.120 1000.000 752.720 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 777.960 1000.000 778.560 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 73.480 1000.000 74.080 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 803.800 1000.000 804.400 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 830.320 1000.000 830.920 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 856.160 1000.000 856.760 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 882.000 1000.000 882.600 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 908.520 1000.000 909.120 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 934.360 1000.000 934.960 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 960.880 1000.000 961.480 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 986.720 1000.000 987.320 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 99.320 1000.000 99.920 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 125.840 1000.000 126.440 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 151.680 1000.000 152.280 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 177.520 1000.000 178.120 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 204.040 1000.000 204.640 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 229.880 1000.000 230.480 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 255.720 1000.000 256.320 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 12.280 1000.000 12.880 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 273.400 1000.000 274.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 299.240 1000.000 299.840 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 325.760 1000.000 326.360 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 351.600 1000.000 352.200 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 378.120 1000.000 378.720 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 403.960 1000.000 404.560 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 429.800 1000.000 430.400 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 456.320 1000.000 456.920 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 482.160 1000.000 482.760 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 508.000 1000.000 508.600 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 38.800 1000.000 39.400 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 534.520 1000.000 535.120 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 560.360 1000.000 560.960 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 586.880 1000.000 587.480 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 612.720 1000.000 613.320 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 638.560 1000.000 639.160 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 665.080 1000.000 665.680 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 690.920 1000.000 691.520 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 716.760 1000.000 717.360 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 743.280 1000.000 743.880 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 769.120 1000.000 769.720 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 64.640 1000.000 65.240 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 795.640 1000.000 796.240 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 821.480 1000.000 822.080 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 847.320 1000.000 847.920 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 873.840 1000.000 874.440 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 899.680 1000.000 900.280 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 925.520 1000.000 926.120 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 952.040 1000.000 952.640 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 977.880 1000.000 978.480 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 90.480 1000.000 91.080 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 117.000 1000.000 117.600 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 142.840 1000.000 143.440 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 169.360 1000.000 169.960 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 195.200 1000.000 195.800 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 221.040 1000.000 221.640 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 247.560 1000.000 248.160 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 995.560 1000.000 996.160 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.230 996.000 993.510 1000.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 0.000 992.130 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 0.000 253.830 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 0.000 361.470 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 0.000 423.110 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 0.000 453.470 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.830 0.000 469.110 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 0.000 669.210 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 0.000 684.390 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 0.000 700.030 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 0.000 730.390 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.750 0.000 746.030 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.930 0.000 761.210 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 0.000 776.850 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.750 0.000 792.030 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.390 0.000 807.670 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.570 0.000 822.850 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.210 0.000 838.490 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 0.000 853.670 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.570 0.000 868.850 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.210 0.000 884.490 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.390 0.000 899.670 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.030 0.000 915.310 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.210 0.000 930.490 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.850 0.000 946.130 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 0.000 530.750 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.030 0.000 961.310 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.670 0.000 976.950 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 0.000 545.930 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 0.000 561.570 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.650 0.000 591.930 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.290 0.000 607.570 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 0.000 622.750 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.110 0.000 638.390 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.720 4.000 664.320 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 679.360 4.000 679.960 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.000 4.000 695.600 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.280 4.000 726.880 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.920 4.000 742.520 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 757.560 4.000 758.160 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.200 4.000 773.800 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 804.480 4.000 805.080 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.960 4.000 523.560 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 820.120 4.000 820.720 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 835.760 4.000 836.360 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 851.400 4.000 852.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 882.680 4.000 883.280 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 898.320 4.000 898.920 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 913.960 4.000 914.560 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 929.600 4.000 930.200 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 960.880 4.000 961.480 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 538.600 4.000 539.200 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 976.520 4.000 977.120 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.160 4.000 992.760 ;
    END
  END la_oenb[31]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 585.520 4.000 586.120 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.160 4.000 601.760 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.800 4.000 617.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.080 4.000 648.680 ;
    END
  END la_oenb[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 996.000 6.810 1000.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 996.000 19.690 1000.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 996.000 72.590 1000.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 996.000 151.250 1000.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 996.000 282.810 1000.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 996.000 296.150 1000.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 996.000 309.030 1000.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 996.000 322.370 1000.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 996.000 335.710 1000.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 996.000 348.590 1000.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 996.000 361.930 1000.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 996.000 374.810 1000.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 996.000 388.150 1000.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 996.000 401.490 1000.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 996.000 164.590 1000.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 996.000 414.370 1000.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 996.000 427.710 1000.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 996.000 440.590 1000.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 996.000 453.930 1000.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 996.000 467.270 1000.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 996.000 480.150 1000.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 996.000 493.490 1000.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 996.000 506.830 1000.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 996.000 519.710 1000.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 996.000 533.050 1000.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 996.000 177.470 1000.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 996.000 545.930 1000.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 996.000 559.270 1000.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 996.000 190.810 1000.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 996.000 204.150 1000.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 996.000 217.030 1000.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 996.000 230.370 1000.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 996.000 243.250 1000.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 996.000 256.590 1000.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 996.000 269.930 1000.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 996.000 45.910 1000.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 996.000 572.610 1000.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 996.000 704.170 1000.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 996.000 717.050 1000.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 996.000 730.390 1000.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.990 996.000 743.270 1000.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.330 996.000 756.610 1000.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 996.000 769.950 1000.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 996.000 782.830 1000.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 996.000 796.170 1000.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.770 996.000 809.050 1000.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 996.000 822.390 1000.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 996.000 585.490 1000.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.450 996.000 835.730 1000.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.330 996.000 848.610 1000.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.670 996.000 861.950 1000.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.550 996.000 874.830 1000.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.890 996.000 888.170 1000.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.230 996.000 901.510 1000.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.110 996.000 914.390 1000.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 996.000 927.730 1000.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 996.000 940.610 1000.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.670 996.000 953.950 1000.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 996.000 598.830 1000.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.010 996.000 967.290 1000.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.890 996.000 980.170 1000.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 996.000 611.710 1000.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 996.000 625.050 1000.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.110 996.000 638.390 1000.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.990 996.000 651.270 1000.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 996.000 664.610 1000.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.210 996.000 677.490 1000.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.550 996.000 690.830 1000.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.160 4.000 210.760 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.720 4.000 273.320 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.000 4.000 304.600 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.280 4.000 335.880 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.560 4.000 367.160 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.120 4.000 429.720 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 460.400 4.000 461.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.680 4.000 492.280 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 4.000 116.920 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 996.000 98.810 1000.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 996.000 111.690 1000.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 996.000 125.030 1000.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 996.000 138.370 1000.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 996.000 33.030 1000.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 996.000 59.250 1000.000 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 987.600 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 987.600 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 987.600 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 987.600 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 987.600 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 987.600 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 987.600 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 987.600 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 987.600 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 987.600 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 987.600 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 987.600 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 987.600 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 945.940 10.880 947.540 987.360 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 792.340 10.880 793.940 987.360 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.740 10.880 640.340 987.360 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 987.360 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 987.360 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 987.360 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 987.360 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 869.140 10.880 870.740 987.360 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 715.540 10.880 717.140 987.360 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.940 10.880 563.540 987.360 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 987.360 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 987.360 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 987.360 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 949.240 10.880 950.840 987.360 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 795.640 10.880 797.240 987.360 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 642.040 10.880 643.640 987.360 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 488.440 10.880 490.040 987.360 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 987.360 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 987.360 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 987.360 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 872.440 10.880 874.040 987.360 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 718.840 10.880 720.440 987.360 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 565.240 10.880 566.840 987.360 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.640 10.880 413.240 987.360 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 987.360 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 987.360 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 952.540 10.880 954.140 987.360 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 798.940 10.880 800.540 987.360 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 645.340 10.880 646.940 987.360 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 491.740 10.880 493.340 987.360 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 987.360 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 987.360 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 987.360 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 875.740 10.880 877.340 987.360 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 722.140 10.880 723.740 987.360 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 568.540 10.880 570.140 987.360 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 414.940 10.880 416.540 987.360 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 987.360 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 987.360 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 994.835 992.035 ;
      LAYER met1 ;
        RECT 5.520 9.560 994.910 997.860 ;
      LAYER met2 ;
        RECT 7.090 995.720 19.130 997.890 ;
        RECT 19.970 995.720 32.470 997.890 ;
        RECT 33.310 995.720 45.350 997.890 ;
        RECT 46.190 995.720 58.690 997.890 ;
        RECT 59.530 995.720 72.030 997.890 ;
        RECT 72.870 995.720 84.910 997.890 ;
        RECT 85.750 995.720 98.250 997.890 ;
        RECT 99.090 995.720 111.130 997.890 ;
        RECT 111.970 995.720 124.470 997.890 ;
        RECT 125.310 995.720 137.810 997.890 ;
        RECT 138.650 995.720 150.690 997.890 ;
        RECT 151.530 995.720 164.030 997.890 ;
        RECT 164.870 995.720 176.910 997.890 ;
        RECT 177.750 995.720 190.250 997.890 ;
        RECT 191.090 995.720 203.590 997.890 ;
        RECT 204.430 995.720 216.470 997.890 ;
        RECT 217.310 995.720 229.810 997.890 ;
        RECT 230.650 995.720 242.690 997.890 ;
        RECT 243.530 995.720 256.030 997.890 ;
        RECT 256.870 995.720 269.370 997.890 ;
        RECT 270.210 995.720 282.250 997.890 ;
        RECT 283.090 995.720 295.590 997.890 ;
        RECT 296.430 995.720 308.470 997.890 ;
        RECT 309.310 995.720 321.810 997.890 ;
        RECT 322.650 995.720 335.150 997.890 ;
        RECT 335.990 995.720 348.030 997.890 ;
        RECT 348.870 995.720 361.370 997.890 ;
        RECT 362.210 995.720 374.250 997.890 ;
        RECT 375.090 995.720 387.590 997.890 ;
        RECT 388.430 995.720 400.930 997.890 ;
        RECT 401.770 995.720 413.810 997.890 ;
        RECT 414.650 995.720 427.150 997.890 ;
        RECT 427.990 995.720 440.030 997.890 ;
        RECT 440.870 995.720 453.370 997.890 ;
        RECT 454.210 995.720 466.710 997.890 ;
        RECT 467.550 995.720 479.590 997.890 ;
        RECT 480.430 995.720 492.930 997.890 ;
        RECT 493.770 995.720 506.270 997.890 ;
        RECT 507.110 995.720 519.150 997.890 ;
        RECT 519.990 995.720 532.490 997.890 ;
        RECT 533.330 995.720 545.370 997.890 ;
        RECT 546.210 995.720 558.710 997.890 ;
        RECT 559.550 995.720 572.050 997.890 ;
        RECT 572.890 995.720 584.930 997.890 ;
        RECT 585.770 995.720 598.270 997.890 ;
        RECT 599.110 995.720 611.150 997.890 ;
        RECT 611.990 995.720 624.490 997.890 ;
        RECT 625.330 995.720 637.830 997.890 ;
        RECT 638.670 995.720 650.710 997.890 ;
        RECT 651.550 995.720 664.050 997.890 ;
        RECT 664.890 995.720 676.930 997.890 ;
        RECT 677.770 995.720 690.270 997.890 ;
        RECT 691.110 995.720 703.610 997.890 ;
        RECT 704.450 995.720 716.490 997.890 ;
        RECT 717.330 995.720 729.830 997.890 ;
        RECT 730.670 995.720 742.710 997.890 ;
        RECT 743.550 995.720 756.050 997.890 ;
        RECT 756.890 995.720 769.390 997.890 ;
        RECT 770.230 995.720 782.270 997.890 ;
        RECT 783.110 995.720 795.610 997.890 ;
        RECT 796.450 995.720 808.490 997.890 ;
        RECT 809.330 995.720 821.830 997.890 ;
        RECT 822.670 995.720 835.170 997.890 ;
        RECT 836.010 995.720 848.050 997.890 ;
        RECT 848.890 995.720 861.390 997.890 ;
        RECT 862.230 995.720 874.270 997.890 ;
        RECT 875.110 995.720 887.610 997.890 ;
        RECT 888.450 995.720 900.950 997.890 ;
        RECT 901.790 995.720 913.830 997.890 ;
        RECT 914.670 995.720 927.170 997.890 ;
        RECT 928.010 995.720 940.050 997.890 ;
        RECT 940.890 995.720 953.390 997.890 ;
        RECT 954.230 995.720 966.730 997.890 ;
        RECT 967.570 995.720 979.610 997.890 ;
        RECT 980.450 995.720 992.950 997.890 ;
        RECT 993.790 995.720 994.890 997.890 ;
        RECT 6.540 4.280 994.890 995.720 ;
        RECT 6.540 4.000 7.170 4.280 ;
        RECT 8.010 4.000 22.350 4.280 ;
        RECT 23.190 4.000 37.530 4.280 ;
        RECT 38.370 4.000 53.170 4.280 ;
        RECT 54.010 4.000 68.350 4.280 ;
        RECT 69.190 4.000 83.990 4.280 ;
        RECT 84.830 4.000 99.170 4.280 ;
        RECT 100.010 4.000 114.810 4.280 ;
        RECT 115.650 4.000 129.990 4.280 ;
        RECT 130.830 4.000 145.630 4.280 ;
        RECT 146.470 4.000 160.810 4.280 ;
        RECT 161.650 4.000 175.990 4.280 ;
        RECT 176.830 4.000 191.630 4.280 ;
        RECT 192.470 4.000 206.810 4.280 ;
        RECT 207.650 4.000 222.450 4.280 ;
        RECT 223.290 4.000 237.630 4.280 ;
        RECT 238.470 4.000 253.270 4.280 ;
        RECT 254.110 4.000 268.450 4.280 ;
        RECT 269.290 4.000 284.090 4.280 ;
        RECT 284.930 4.000 299.270 4.280 ;
        RECT 300.110 4.000 314.450 4.280 ;
        RECT 315.290 4.000 330.090 4.280 ;
        RECT 330.930 4.000 345.270 4.280 ;
        RECT 346.110 4.000 360.910 4.280 ;
        RECT 361.750 4.000 376.090 4.280 ;
        RECT 376.930 4.000 391.730 4.280 ;
        RECT 392.570 4.000 406.910 4.280 ;
        RECT 407.750 4.000 422.550 4.280 ;
        RECT 423.390 4.000 437.730 4.280 ;
        RECT 438.570 4.000 452.910 4.280 ;
        RECT 453.750 4.000 468.550 4.280 ;
        RECT 469.390 4.000 483.730 4.280 ;
        RECT 484.570 4.000 499.370 4.280 ;
        RECT 500.210 4.000 514.550 4.280 ;
        RECT 515.390 4.000 530.190 4.280 ;
        RECT 531.030 4.000 545.370 4.280 ;
        RECT 546.210 4.000 561.010 4.280 ;
        RECT 561.850 4.000 576.190 4.280 ;
        RECT 577.030 4.000 591.370 4.280 ;
        RECT 592.210 4.000 607.010 4.280 ;
        RECT 607.850 4.000 622.190 4.280 ;
        RECT 623.030 4.000 637.830 4.280 ;
        RECT 638.670 4.000 653.010 4.280 ;
        RECT 653.850 4.000 668.650 4.280 ;
        RECT 669.490 4.000 683.830 4.280 ;
        RECT 684.670 4.000 699.470 4.280 ;
        RECT 700.310 4.000 714.650 4.280 ;
        RECT 715.490 4.000 729.830 4.280 ;
        RECT 730.670 4.000 745.470 4.280 ;
        RECT 746.310 4.000 760.650 4.280 ;
        RECT 761.490 4.000 776.290 4.280 ;
        RECT 777.130 4.000 791.470 4.280 ;
        RECT 792.310 4.000 807.110 4.280 ;
        RECT 807.950 4.000 822.290 4.280 ;
        RECT 823.130 4.000 837.930 4.280 ;
        RECT 838.770 4.000 853.110 4.280 ;
        RECT 853.950 4.000 868.290 4.280 ;
        RECT 869.130 4.000 883.930 4.280 ;
        RECT 884.770 4.000 899.110 4.280 ;
        RECT 899.950 4.000 914.750 4.280 ;
        RECT 915.590 4.000 929.930 4.280 ;
        RECT 930.770 4.000 945.570 4.280 ;
        RECT 946.410 4.000 960.750 4.280 ;
        RECT 961.590 4.000 976.390 4.280 ;
        RECT 977.230 4.000 991.570 4.280 ;
        RECT 992.410 4.000 994.890 4.280 ;
      LAYER met3 ;
        RECT 4.000 995.160 995.600 996.025 ;
        RECT 4.000 993.160 996.000 995.160 ;
        RECT 4.400 991.760 996.000 993.160 ;
        RECT 4.000 987.720 996.000 991.760 ;
        RECT 4.000 986.320 995.600 987.720 ;
        RECT 4.000 978.880 996.000 986.320 ;
        RECT 4.000 977.520 995.600 978.880 ;
        RECT 4.400 977.480 995.600 977.520 ;
        RECT 4.400 976.120 996.000 977.480 ;
        RECT 4.000 970.040 996.000 976.120 ;
        RECT 4.000 968.640 995.600 970.040 ;
        RECT 4.000 961.880 996.000 968.640 ;
        RECT 4.400 960.480 995.600 961.880 ;
        RECT 4.000 953.040 996.000 960.480 ;
        RECT 4.000 951.640 995.600 953.040 ;
        RECT 4.000 946.240 996.000 951.640 ;
        RECT 4.400 944.840 996.000 946.240 ;
        RECT 4.000 944.200 996.000 944.840 ;
        RECT 4.000 942.800 995.600 944.200 ;
        RECT 4.000 935.360 996.000 942.800 ;
        RECT 4.000 933.960 995.600 935.360 ;
        RECT 4.000 930.600 996.000 933.960 ;
        RECT 4.400 929.200 996.000 930.600 ;
        RECT 4.000 926.520 996.000 929.200 ;
        RECT 4.000 925.120 995.600 926.520 ;
        RECT 4.000 918.360 996.000 925.120 ;
        RECT 4.000 916.960 995.600 918.360 ;
        RECT 4.000 914.960 996.000 916.960 ;
        RECT 4.400 913.560 996.000 914.960 ;
        RECT 4.000 909.520 996.000 913.560 ;
        RECT 4.000 908.120 995.600 909.520 ;
        RECT 4.000 900.680 996.000 908.120 ;
        RECT 4.000 899.320 995.600 900.680 ;
        RECT 4.400 899.280 995.600 899.320 ;
        RECT 4.400 897.920 996.000 899.280 ;
        RECT 4.000 891.840 996.000 897.920 ;
        RECT 4.000 890.440 995.600 891.840 ;
        RECT 4.000 883.680 996.000 890.440 ;
        RECT 4.400 883.000 996.000 883.680 ;
        RECT 4.400 882.280 995.600 883.000 ;
        RECT 4.000 881.600 995.600 882.280 ;
        RECT 4.000 874.840 996.000 881.600 ;
        RECT 4.000 873.440 995.600 874.840 ;
        RECT 4.000 868.040 996.000 873.440 ;
        RECT 4.400 866.640 996.000 868.040 ;
        RECT 4.000 866.000 996.000 866.640 ;
        RECT 4.000 864.600 995.600 866.000 ;
        RECT 4.000 857.160 996.000 864.600 ;
        RECT 4.000 855.760 995.600 857.160 ;
        RECT 4.000 852.400 996.000 855.760 ;
        RECT 4.400 851.000 996.000 852.400 ;
        RECT 4.000 848.320 996.000 851.000 ;
        RECT 4.000 846.920 995.600 848.320 ;
        RECT 4.000 839.480 996.000 846.920 ;
        RECT 4.000 838.080 995.600 839.480 ;
        RECT 4.000 836.760 996.000 838.080 ;
        RECT 4.400 835.360 996.000 836.760 ;
        RECT 4.000 831.320 996.000 835.360 ;
        RECT 4.000 829.920 995.600 831.320 ;
        RECT 4.000 822.480 996.000 829.920 ;
        RECT 4.000 821.120 995.600 822.480 ;
        RECT 4.400 821.080 995.600 821.120 ;
        RECT 4.400 819.720 996.000 821.080 ;
        RECT 4.000 813.640 996.000 819.720 ;
        RECT 4.000 812.240 995.600 813.640 ;
        RECT 4.000 805.480 996.000 812.240 ;
        RECT 4.400 804.800 996.000 805.480 ;
        RECT 4.400 804.080 995.600 804.800 ;
        RECT 4.000 803.400 995.600 804.080 ;
        RECT 4.000 796.640 996.000 803.400 ;
        RECT 4.000 795.240 995.600 796.640 ;
        RECT 4.000 789.840 996.000 795.240 ;
        RECT 4.400 788.440 996.000 789.840 ;
        RECT 4.000 787.800 996.000 788.440 ;
        RECT 4.000 786.400 995.600 787.800 ;
        RECT 4.000 778.960 996.000 786.400 ;
        RECT 4.000 777.560 995.600 778.960 ;
        RECT 4.000 774.200 996.000 777.560 ;
        RECT 4.400 772.800 996.000 774.200 ;
        RECT 4.000 770.120 996.000 772.800 ;
        RECT 4.000 768.720 995.600 770.120 ;
        RECT 4.000 761.280 996.000 768.720 ;
        RECT 4.000 759.880 995.600 761.280 ;
        RECT 4.000 758.560 996.000 759.880 ;
        RECT 4.400 757.160 996.000 758.560 ;
        RECT 4.000 753.120 996.000 757.160 ;
        RECT 4.000 751.720 995.600 753.120 ;
        RECT 4.000 744.280 996.000 751.720 ;
        RECT 4.000 742.920 995.600 744.280 ;
        RECT 4.400 742.880 995.600 742.920 ;
        RECT 4.400 741.520 996.000 742.880 ;
        RECT 4.000 735.440 996.000 741.520 ;
        RECT 4.000 734.040 995.600 735.440 ;
        RECT 4.000 727.280 996.000 734.040 ;
        RECT 4.400 726.600 996.000 727.280 ;
        RECT 4.400 725.880 995.600 726.600 ;
        RECT 4.000 725.200 995.600 725.880 ;
        RECT 4.000 717.760 996.000 725.200 ;
        RECT 4.000 716.360 995.600 717.760 ;
        RECT 4.000 711.640 996.000 716.360 ;
        RECT 4.400 710.240 996.000 711.640 ;
        RECT 4.000 709.600 996.000 710.240 ;
        RECT 4.000 708.200 995.600 709.600 ;
        RECT 4.000 700.760 996.000 708.200 ;
        RECT 4.000 699.360 995.600 700.760 ;
        RECT 4.000 696.000 996.000 699.360 ;
        RECT 4.400 694.600 996.000 696.000 ;
        RECT 4.000 691.920 996.000 694.600 ;
        RECT 4.000 690.520 995.600 691.920 ;
        RECT 4.000 683.080 996.000 690.520 ;
        RECT 4.000 681.680 995.600 683.080 ;
        RECT 4.000 680.360 996.000 681.680 ;
        RECT 4.400 678.960 996.000 680.360 ;
        RECT 4.000 674.240 996.000 678.960 ;
        RECT 4.000 672.840 995.600 674.240 ;
        RECT 4.000 666.080 996.000 672.840 ;
        RECT 4.000 664.720 995.600 666.080 ;
        RECT 4.400 664.680 995.600 664.720 ;
        RECT 4.400 663.320 996.000 664.680 ;
        RECT 4.000 657.240 996.000 663.320 ;
        RECT 4.000 655.840 995.600 657.240 ;
        RECT 4.000 649.080 996.000 655.840 ;
        RECT 4.400 648.400 996.000 649.080 ;
        RECT 4.400 647.680 995.600 648.400 ;
        RECT 4.000 647.000 995.600 647.680 ;
        RECT 4.000 639.560 996.000 647.000 ;
        RECT 4.000 638.160 995.600 639.560 ;
        RECT 4.000 633.440 996.000 638.160 ;
        RECT 4.400 632.040 996.000 633.440 ;
        RECT 4.000 630.720 996.000 632.040 ;
        RECT 4.000 629.320 995.600 630.720 ;
        RECT 4.000 622.560 996.000 629.320 ;
        RECT 4.000 621.160 995.600 622.560 ;
        RECT 4.000 617.800 996.000 621.160 ;
        RECT 4.400 616.400 996.000 617.800 ;
        RECT 4.000 613.720 996.000 616.400 ;
        RECT 4.000 612.320 995.600 613.720 ;
        RECT 4.000 604.880 996.000 612.320 ;
        RECT 4.000 603.480 995.600 604.880 ;
        RECT 4.000 602.160 996.000 603.480 ;
        RECT 4.400 600.760 996.000 602.160 ;
        RECT 4.000 596.040 996.000 600.760 ;
        RECT 4.000 594.640 995.600 596.040 ;
        RECT 4.000 587.880 996.000 594.640 ;
        RECT 4.000 586.520 995.600 587.880 ;
        RECT 4.400 586.480 995.600 586.520 ;
        RECT 4.400 585.120 996.000 586.480 ;
        RECT 4.000 579.040 996.000 585.120 ;
        RECT 4.000 577.640 995.600 579.040 ;
        RECT 4.000 570.880 996.000 577.640 ;
        RECT 4.400 570.200 996.000 570.880 ;
        RECT 4.400 569.480 995.600 570.200 ;
        RECT 4.000 568.800 995.600 569.480 ;
        RECT 4.000 561.360 996.000 568.800 ;
        RECT 4.000 559.960 995.600 561.360 ;
        RECT 4.000 555.240 996.000 559.960 ;
        RECT 4.400 553.840 996.000 555.240 ;
        RECT 4.000 552.520 996.000 553.840 ;
        RECT 4.000 551.120 995.600 552.520 ;
        RECT 4.000 544.360 996.000 551.120 ;
        RECT 4.000 542.960 995.600 544.360 ;
        RECT 4.000 539.600 996.000 542.960 ;
        RECT 4.400 538.200 996.000 539.600 ;
        RECT 4.000 535.520 996.000 538.200 ;
        RECT 4.000 534.120 995.600 535.520 ;
        RECT 4.000 526.680 996.000 534.120 ;
        RECT 4.000 525.280 995.600 526.680 ;
        RECT 4.000 523.960 996.000 525.280 ;
        RECT 4.400 522.560 996.000 523.960 ;
        RECT 4.000 517.840 996.000 522.560 ;
        RECT 4.000 516.440 995.600 517.840 ;
        RECT 4.000 509.000 996.000 516.440 ;
        RECT 4.000 508.320 995.600 509.000 ;
        RECT 4.400 507.600 995.600 508.320 ;
        RECT 4.400 506.920 996.000 507.600 ;
        RECT 4.000 500.840 996.000 506.920 ;
        RECT 4.000 499.440 995.600 500.840 ;
        RECT 4.000 492.680 996.000 499.440 ;
        RECT 4.400 492.000 996.000 492.680 ;
        RECT 4.400 491.280 995.600 492.000 ;
        RECT 4.000 490.600 995.600 491.280 ;
        RECT 4.000 483.160 996.000 490.600 ;
        RECT 4.000 481.760 995.600 483.160 ;
        RECT 4.000 477.040 996.000 481.760 ;
        RECT 4.400 475.640 996.000 477.040 ;
        RECT 4.000 474.320 996.000 475.640 ;
        RECT 4.000 472.920 995.600 474.320 ;
        RECT 4.000 465.480 996.000 472.920 ;
        RECT 4.000 464.080 995.600 465.480 ;
        RECT 4.000 461.400 996.000 464.080 ;
        RECT 4.400 460.000 996.000 461.400 ;
        RECT 4.000 457.320 996.000 460.000 ;
        RECT 4.000 455.920 995.600 457.320 ;
        RECT 4.000 448.480 996.000 455.920 ;
        RECT 4.000 447.080 995.600 448.480 ;
        RECT 4.000 445.760 996.000 447.080 ;
        RECT 4.400 444.360 996.000 445.760 ;
        RECT 4.000 439.640 996.000 444.360 ;
        RECT 4.000 438.240 995.600 439.640 ;
        RECT 4.000 430.800 996.000 438.240 ;
        RECT 4.000 430.120 995.600 430.800 ;
        RECT 4.400 429.400 995.600 430.120 ;
        RECT 4.400 428.720 996.000 429.400 ;
        RECT 4.000 421.960 996.000 428.720 ;
        RECT 4.000 420.560 995.600 421.960 ;
        RECT 4.000 414.480 996.000 420.560 ;
        RECT 4.400 413.800 996.000 414.480 ;
        RECT 4.400 413.080 995.600 413.800 ;
        RECT 4.000 412.400 995.600 413.080 ;
        RECT 4.000 404.960 996.000 412.400 ;
        RECT 4.000 403.560 995.600 404.960 ;
        RECT 4.000 398.840 996.000 403.560 ;
        RECT 4.400 397.440 996.000 398.840 ;
        RECT 4.000 396.120 996.000 397.440 ;
        RECT 4.000 394.720 995.600 396.120 ;
        RECT 4.000 387.280 996.000 394.720 ;
        RECT 4.000 385.880 995.600 387.280 ;
        RECT 4.000 383.200 996.000 385.880 ;
        RECT 4.400 381.800 996.000 383.200 ;
        RECT 4.000 379.120 996.000 381.800 ;
        RECT 4.000 377.720 995.600 379.120 ;
        RECT 4.000 370.280 996.000 377.720 ;
        RECT 4.000 368.880 995.600 370.280 ;
        RECT 4.000 367.560 996.000 368.880 ;
        RECT 4.400 366.160 996.000 367.560 ;
        RECT 4.000 361.440 996.000 366.160 ;
        RECT 4.000 360.040 995.600 361.440 ;
        RECT 4.000 352.600 996.000 360.040 ;
        RECT 4.000 351.920 995.600 352.600 ;
        RECT 4.400 351.200 995.600 351.920 ;
        RECT 4.400 350.520 996.000 351.200 ;
        RECT 4.000 343.760 996.000 350.520 ;
        RECT 4.000 342.360 995.600 343.760 ;
        RECT 4.000 336.280 996.000 342.360 ;
        RECT 4.400 335.600 996.000 336.280 ;
        RECT 4.400 334.880 995.600 335.600 ;
        RECT 4.000 334.200 995.600 334.880 ;
        RECT 4.000 326.760 996.000 334.200 ;
        RECT 4.000 325.360 995.600 326.760 ;
        RECT 4.000 320.640 996.000 325.360 ;
        RECT 4.400 319.240 996.000 320.640 ;
        RECT 4.000 317.920 996.000 319.240 ;
        RECT 4.000 316.520 995.600 317.920 ;
        RECT 4.000 309.080 996.000 316.520 ;
        RECT 4.000 307.680 995.600 309.080 ;
        RECT 4.000 305.000 996.000 307.680 ;
        RECT 4.400 303.600 996.000 305.000 ;
        RECT 4.000 300.240 996.000 303.600 ;
        RECT 4.000 298.840 995.600 300.240 ;
        RECT 4.000 292.080 996.000 298.840 ;
        RECT 4.000 290.680 995.600 292.080 ;
        RECT 4.000 289.360 996.000 290.680 ;
        RECT 4.400 287.960 996.000 289.360 ;
        RECT 4.000 283.240 996.000 287.960 ;
        RECT 4.000 281.840 995.600 283.240 ;
        RECT 4.000 274.400 996.000 281.840 ;
        RECT 4.000 273.720 995.600 274.400 ;
        RECT 4.400 273.000 995.600 273.720 ;
        RECT 4.400 272.320 996.000 273.000 ;
        RECT 4.000 265.560 996.000 272.320 ;
        RECT 4.000 264.160 995.600 265.560 ;
        RECT 4.000 258.080 996.000 264.160 ;
        RECT 4.400 256.720 996.000 258.080 ;
        RECT 4.400 256.680 995.600 256.720 ;
        RECT 4.000 255.320 995.600 256.680 ;
        RECT 4.000 248.560 996.000 255.320 ;
        RECT 4.000 247.160 995.600 248.560 ;
        RECT 4.000 242.440 996.000 247.160 ;
        RECT 4.400 241.040 996.000 242.440 ;
        RECT 4.000 239.720 996.000 241.040 ;
        RECT 4.000 238.320 995.600 239.720 ;
        RECT 4.000 230.880 996.000 238.320 ;
        RECT 4.000 229.480 995.600 230.880 ;
        RECT 4.000 226.800 996.000 229.480 ;
        RECT 4.400 225.400 996.000 226.800 ;
        RECT 4.000 222.040 996.000 225.400 ;
        RECT 4.000 220.640 995.600 222.040 ;
        RECT 4.000 213.200 996.000 220.640 ;
        RECT 4.000 211.800 995.600 213.200 ;
        RECT 4.000 211.160 996.000 211.800 ;
        RECT 4.400 209.760 996.000 211.160 ;
        RECT 4.000 205.040 996.000 209.760 ;
        RECT 4.000 203.640 995.600 205.040 ;
        RECT 4.000 196.200 996.000 203.640 ;
        RECT 4.000 195.520 995.600 196.200 ;
        RECT 4.400 194.800 995.600 195.520 ;
        RECT 4.400 194.120 996.000 194.800 ;
        RECT 4.000 187.360 996.000 194.120 ;
        RECT 4.000 185.960 995.600 187.360 ;
        RECT 4.000 179.880 996.000 185.960 ;
        RECT 4.400 178.520 996.000 179.880 ;
        RECT 4.400 178.480 995.600 178.520 ;
        RECT 4.000 177.120 995.600 178.480 ;
        RECT 4.000 170.360 996.000 177.120 ;
        RECT 4.000 168.960 995.600 170.360 ;
        RECT 4.000 164.240 996.000 168.960 ;
        RECT 4.400 162.840 996.000 164.240 ;
        RECT 4.000 161.520 996.000 162.840 ;
        RECT 4.000 160.120 995.600 161.520 ;
        RECT 4.000 152.680 996.000 160.120 ;
        RECT 4.000 151.280 995.600 152.680 ;
        RECT 4.000 148.600 996.000 151.280 ;
        RECT 4.400 147.200 996.000 148.600 ;
        RECT 4.000 143.840 996.000 147.200 ;
        RECT 4.000 142.440 995.600 143.840 ;
        RECT 4.000 135.000 996.000 142.440 ;
        RECT 4.000 133.600 995.600 135.000 ;
        RECT 4.000 132.960 996.000 133.600 ;
        RECT 4.400 131.560 996.000 132.960 ;
        RECT 4.000 126.840 996.000 131.560 ;
        RECT 4.000 125.440 995.600 126.840 ;
        RECT 4.000 118.000 996.000 125.440 ;
        RECT 4.000 117.320 995.600 118.000 ;
        RECT 4.400 116.600 995.600 117.320 ;
        RECT 4.400 115.920 996.000 116.600 ;
        RECT 4.000 109.160 996.000 115.920 ;
        RECT 4.000 107.760 995.600 109.160 ;
        RECT 4.000 101.680 996.000 107.760 ;
        RECT 4.400 100.320 996.000 101.680 ;
        RECT 4.400 100.280 995.600 100.320 ;
        RECT 4.000 98.920 995.600 100.280 ;
        RECT 4.000 91.480 996.000 98.920 ;
        RECT 4.000 90.080 995.600 91.480 ;
        RECT 4.000 86.040 996.000 90.080 ;
        RECT 4.400 84.640 996.000 86.040 ;
        RECT 4.000 83.320 996.000 84.640 ;
        RECT 4.000 81.920 995.600 83.320 ;
        RECT 4.000 74.480 996.000 81.920 ;
        RECT 4.000 73.080 995.600 74.480 ;
        RECT 4.000 70.400 996.000 73.080 ;
        RECT 4.400 69.000 996.000 70.400 ;
        RECT 4.000 65.640 996.000 69.000 ;
        RECT 4.000 64.240 995.600 65.640 ;
        RECT 4.000 56.800 996.000 64.240 ;
        RECT 4.000 55.400 995.600 56.800 ;
        RECT 4.000 54.760 996.000 55.400 ;
        RECT 4.400 53.360 996.000 54.760 ;
        RECT 4.000 47.960 996.000 53.360 ;
        RECT 4.000 46.560 995.600 47.960 ;
        RECT 4.000 39.800 996.000 46.560 ;
        RECT 4.000 39.120 995.600 39.800 ;
        RECT 4.400 38.400 995.600 39.120 ;
        RECT 4.400 37.720 996.000 38.400 ;
        RECT 4.000 30.960 996.000 37.720 ;
        RECT 4.000 29.560 995.600 30.960 ;
        RECT 4.000 23.480 996.000 29.560 ;
        RECT 4.400 22.120 996.000 23.480 ;
        RECT 4.400 22.080 995.600 22.120 ;
        RECT 4.000 20.720 995.600 22.080 ;
        RECT 4.000 13.280 996.000 20.720 ;
        RECT 4.000 11.880 995.600 13.280 ;
        RECT 4.000 8.520 996.000 11.880 ;
        RECT 4.400 7.120 996.000 8.520 ;
        RECT 4.000 5.120 996.000 7.120 ;
        RECT 4.000 4.255 995.600 5.120 ;
      LAYER met4 ;
        RECT 157.615 123.935 174.240 966.105 ;
        RECT 176.640 123.935 177.540 966.105 ;
        RECT 179.940 123.935 180.840 966.105 ;
        RECT 183.240 123.935 184.140 966.105 ;
        RECT 186.540 123.935 251.040 966.105 ;
        RECT 253.440 123.935 254.340 966.105 ;
        RECT 256.740 123.935 257.640 966.105 ;
        RECT 260.040 123.935 260.940 966.105 ;
        RECT 263.340 123.935 327.840 966.105 ;
        RECT 330.240 123.935 331.140 966.105 ;
        RECT 333.540 123.935 334.440 966.105 ;
        RECT 336.840 123.935 337.740 966.105 ;
        RECT 340.140 123.935 404.640 966.105 ;
        RECT 407.040 123.935 407.940 966.105 ;
        RECT 410.340 123.935 411.240 966.105 ;
        RECT 413.640 123.935 414.540 966.105 ;
        RECT 416.940 123.935 481.440 966.105 ;
        RECT 483.840 123.935 484.740 966.105 ;
        RECT 487.140 123.935 488.040 966.105 ;
        RECT 490.440 123.935 491.340 966.105 ;
        RECT 493.740 123.935 558.240 966.105 ;
        RECT 560.640 123.935 561.540 966.105 ;
        RECT 563.940 123.935 564.840 966.105 ;
        RECT 567.240 123.935 568.140 966.105 ;
        RECT 570.540 123.935 635.040 966.105 ;
        RECT 637.440 123.935 638.340 966.105 ;
        RECT 640.740 123.935 641.640 966.105 ;
        RECT 644.040 123.935 644.940 966.105 ;
        RECT 647.340 123.935 711.840 966.105 ;
        RECT 714.240 123.935 715.140 966.105 ;
        RECT 717.540 123.935 718.440 966.105 ;
        RECT 720.840 123.935 721.740 966.105 ;
        RECT 724.140 123.935 788.640 966.105 ;
        RECT 791.040 123.935 791.940 966.105 ;
        RECT 794.340 123.935 795.240 966.105 ;
        RECT 797.640 123.935 798.540 966.105 ;
        RECT 800.940 123.935 865.440 966.105 ;
        RECT 867.840 123.935 868.740 966.105 ;
        RECT 871.140 123.935 872.040 966.105 ;
        RECT 874.440 123.935 875.340 966.105 ;
        RECT 877.740 123.935 892.105 966.105 ;
  END
END wrapper_sha1
END LIBRARY

