VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapper_sha1
  CLASS BLOCK ;
  FOREIGN wrapper_sha1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 800.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 796.000 69.370 800.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 3.440 800.000 4.040 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 211.520 800.000 212.120 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 232.600 800.000 233.200 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 253.680 800.000 254.280 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 274.080 800.000 274.680 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 295.160 800.000 295.760 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 316.240 800.000 316.840 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 336.640 800.000 337.240 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 357.720 800.000 358.320 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 378.800 800.000 379.400 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 399.200 800.000 399.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 23.840 800.000 24.440 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 420.280 800.000 420.880 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 441.360 800.000 441.960 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 461.760 800.000 462.360 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 482.840 800.000 483.440 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 503.920 800.000 504.520 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 524.320 800.000 524.920 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 545.400 800.000 546.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 566.480 800.000 567.080 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 586.880 800.000 587.480 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 607.960 800.000 608.560 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 44.920 800.000 45.520 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 629.040 800.000 629.640 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 650.120 800.000 650.720 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 670.520 800.000 671.120 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 691.600 800.000 692.200 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 712.680 800.000 713.280 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 733.080 800.000 733.680 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 754.160 800.000 754.760 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 775.240 800.000 775.840 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 66.000 800.000 66.600 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 86.400 800.000 87.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 107.480 800.000 108.080 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 128.560 800.000 129.160 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 148.960 800.000 149.560 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 170.040 800.000 170.640 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 191.120 800.000 191.720 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 17.040 800.000 17.640 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 225.800 800.000 226.400 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 246.200 800.000 246.800 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 267.280 800.000 267.880 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 288.360 800.000 288.960 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 308.760 800.000 309.360 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 329.840 800.000 330.440 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 350.920 800.000 351.520 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 371.320 800.000 371.920 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 392.400 800.000 393.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 413.480 800.000 414.080 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 38.120 800.000 38.720 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 434.560 800.000 435.160 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 454.960 800.000 455.560 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 476.040 800.000 476.640 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 497.120 800.000 497.720 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 517.520 800.000 518.120 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 538.600 800.000 539.200 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 559.680 800.000 560.280 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 580.080 800.000 580.680 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 601.160 800.000 601.760 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 622.240 800.000 622.840 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 58.520 800.000 59.120 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 642.640 800.000 643.240 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 663.720 800.000 664.320 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 684.800 800.000 685.400 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 705.200 800.000 705.800 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 726.280 800.000 726.880 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 747.360 800.000 747.960 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 767.760 800.000 768.360 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 788.840 800.000 789.440 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 79.600 800.000 80.200 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 100.680 800.000 101.280 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 121.080 800.000 121.680 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 142.160 800.000 142.760 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 163.240 800.000 163.840 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 183.640 800.000 184.240 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 204.720 800.000 205.320 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 10.240 800.000 10.840 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 219.000 800.000 219.600 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 239.400 800.000 240.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 260.480 800.000 261.080 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 281.560 800.000 282.160 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 301.960 800.000 302.560 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 323.040 800.000 323.640 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 344.120 800.000 344.720 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 364.520 800.000 365.120 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 385.600 800.000 386.200 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 406.680 800.000 407.280 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 30.640 800.000 31.240 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 427.080 800.000 427.680 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 448.160 800.000 448.760 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 469.240 800.000 469.840 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 489.640 800.000 490.240 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 510.720 800.000 511.320 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 531.800 800.000 532.400 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 552.200 800.000 552.800 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 573.280 800.000 573.880 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 594.360 800.000 594.960 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 614.760 800.000 615.360 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 51.720 800.000 52.320 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 635.840 800.000 636.440 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 656.920 800.000 657.520 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 677.320 800.000 677.920 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 698.400 800.000 699.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 719.480 800.000 720.080 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 739.880 800.000 740.480 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 760.960 800.000 761.560 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 782.040 800.000 782.640 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 72.800 800.000 73.400 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 93.200 800.000 93.800 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 114.280 800.000 114.880 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 135.360 800.000 135.960 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 155.760 800.000 156.360 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 176.840 800.000 177.440 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 197.920 800.000 198.520 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.630 0.000 781.910 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 795.640 800.000 796.240 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 0.000 321.450 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 0.000 381.710 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.790 0.000 527.070 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 0.000 539.490 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 0.000 551.450 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 0.000 575.830 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 0.000 587.790 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 0.000 600.210 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 0.000 624.130 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 0.000 636.550 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.230 0.000 648.510 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 0.000 672.890 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.570 0.000 684.850 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.530 0.000 696.810 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 0.000 709.230 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.910 0.000 721.190 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 0.000 733.150 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 0.000 745.570 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.250 0.000 757.530 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.210 0.000 769.490 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 0.000 466.810 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 0.000 503.150 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.000 4.000 406.600 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 543.360 4.000 543.960 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 555.600 4.000 556.200 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.760 4.000 581.360 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.000 4.000 593.600 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.920 4.000 606.520 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.160 4.000 618.760 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 630.400 4.000 631.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.800 4.000 668.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.720 4.000 681.320 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 692.960 4.000 693.560 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 718.120 4.000 718.720 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 730.360 4.000 730.960 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.280 4.000 743.880 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 755.520 4.000 756.120 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 767.760 4.000 768.360 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 430.480 4.000 431.080 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.680 4.000 781.280 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.920 4.000 793.520 ;
    END
  END la_oenb[31]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.800 4.000 481.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.960 4.000 506.560 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END la_oenb[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 796.000 5.430 800.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 796.000 16.010 800.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 796.000 58.330 800.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 796.000 122.730 800.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 796.000 228.990 800.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 796.000 240.030 800.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 796.000 250.610 800.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 796.000 261.190 800.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 796.000 271.770 800.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 796.000 282.350 800.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 796.000 293.390 800.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 796.000 303.970 800.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 796.000 314.550 800.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 796.000 325.130 800.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 796.000 133.310 800.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 796.000 335.710 800.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 796.000 346.290 800.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 796.000 357.330 800.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 796.000 367.910 800.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 796.000 378.490 800.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 796.000 389.070 800.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 796.000 399.650 800.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 796.000 410.690 800.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 796.000 421.270 800.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 796.000 431.850 800.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 796.000 143.890 800.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 796.000 442.430 800.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 796.000 453.010 800.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 796.000 154.470 800.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 796.000 165.050 800.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 796.000 175.630 800.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 796.000 186.670 800.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 796.000 197.250 800.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 796.000 207.830 800.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 796.000 218.410 800.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 796.000 37.170 800.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 796.000 464.050 800.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 796.000 570.310 800.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 796.000 581.350 800.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.650 796.000 591.930 800.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 796.000 602.510 800.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 796.000 613.090 800.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 796.000 623.670 800.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 796.000 634.710 800.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 796.000 645.290 800.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.590 796.000 655.870 800.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.170 796.000 666.450 800.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 796.000 474.630 800.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 796.000 677.030 800.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 796.000 687.610 800.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.370 796.000 698.650 800.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 796.000 709.230 800.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.530 796.000 719.810 800.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 796.000 730.390 800.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 796.000 740.970 800.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.730 796.000 752.010 800.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.310 796.000 762.590 800.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 796.000 773.170 800.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 796.000 485.210 800.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.470 796.000 783.750 800.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 796.000 794.330 800.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 796.000 495.790 800.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 796.000 506.370 800.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 796.000 516.950 800.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 796.000 527.990 800.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 796.000 538.570 800.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.870 796.000 549.150 800.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 796.000 559.730 800.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.320 4.000 218.920 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.560 4.000 231.160 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.680 4.000 356.280 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.920 4.000 368.520 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 796.000 79.950 800.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 796.000 90.530 800.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 796.000 101.110 800.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 796.000 111.690 800.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 796.000 26.590 800.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 796.000 47.750 800.000 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.740 10.880 640.340 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 788.800 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 715.540 10.880 717.140 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.940 10.880 563.540 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 788.800 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 642.040 10.880 643.640 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 488.440 10.880 490.040 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 788.800 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 718.840 10.880 720.440 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 565.240 10.880 566.840 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.640 10.880 413.240 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 788.800 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 645.340 10.880 646.940 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 491.740 10.880 493.340 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 788.800 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 722.140 10.880 723.740 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 568.540 10.880 570.140 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 414.940 10.880 416.540 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 788.800 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 1.065 1.105 795.195 795.175 ;
      LAYER met1 ;
        RECT 0.070 0.040 799.870 795.560 ;
      LAYER met2 ;
        RECT 0.090 795.720 4.870 796.125 ;
        RECT 5.710 795.720 15.450 796.125 ;
        RECT 16.290 795.720 26.030 796.125 ;
        RECT 26.870 795.720 36.610 796.125 ;
        RECT 37.450 795.720 47.190 796.125 ;
        RECT 48.030 795.720 57.770 796.125 ;
        RECT 58.610 795.720 68.810 796.125 ;
        RECT 69.650 795.720 79.390 796.125 ;
        RECT 80.230 795.720 89.970 796.125 ;
        RECT 90.810 795.720 100.550 796.125 ;
        RECT 101.390 795.720 111.130 796.125 ;
        RECT 111.970 795.720 122.170 796.125 ;
        RECT 123.010 795.720 132.750 796.125 ;
        RECT 133.590 795.720 143.330 796.125 ;
        RECT 144.170 795.720 153.910 796.125 ;
        RECT 154.750 795.720 164.490 796.125 ;
        RECT 165.330 795.720 175.070 796.125 ;
        RECT 175.910 795.720 186.110 796.125 ;
        RECT 186.950 795.720 196.690 796.125 ;
        RECT 197.530 795.720 207.270 796.125 ;
        RECT 208.110 795.720 217.850 796.125 ;
        RECT 218.690 795.720 228.430 796.125 ;
        RECT 229.270 795.720 239.470 796.125 ;
        RECT 240.310 795.720 250.050 796.125 ;
        RECT 250.890 795.720 260.630 796.125 ;
        RECT 261.470 795.720 271.210 796.125 ;
        RECT 272.050 795.720 281.790 796.125 ;
        RECT 282.630 795.720 292.830 796.125 ;
        RECT 293.670 795.720 303.410 796.125 ;
        RECT 304.250 795.720 313.990 796.125 ;
        RECT 314.830 795.720 324.570 796.125 ;
        RECT 325.410 795.720 335.150 796.125 ;
        RECT 335.990 795.720 345.730 796.125 ;
        RECT 346.570 795.720 356.770 796.125 ;
        RECT 357.610 795.720 367.350 796.125 ;
        RECT 368.190 795.720 377.930 796.125 ;
        RECT 378.770 795.720 388.510 796.125 ;
        RECT 389.350 795.720 399.090 796.125 ;
        RECT 399.930 795.720 410.130 796.125 ;
        RECT 410.970 795.720 420.710 796.125 ;
        RECT 421.550 795.720 431.290 796.125 ;
        RECT 432.130 795.720 441.870 796.125 ;
        RECT 442.710 795.720 452.450 796.125 ;
        RECT 453.290 795.720 463.490 796.125 ;
        RECT 464.330 795.720 474.070 796.125 ;
        RECT 474.910 795.720 484.650 796.125 ;
        RECT 485.490 795.720 495.230 796.125 ;
        RECT 496.070 795.720 505.810 796.125 ;
        RECT 506.650 795.720 516.390 796.125 ;
        RECT 517.230 795.720 527.430 796.125 ;
        RECT 528.270 795.720 538.010 796.125 ;
        RECT 538.850 795.720 548.590 796.125 ;
        RECT 549.430 795.720 559.170 796.125 ;
        RECT 560.010 795.720 569.750 796.125 ;
        RECT 570.590 795.720 580.790 796.125 ;
        RECT 581.630 795.720 591.370 796.125 ;
        RECT 592.210 795.720 601.950 796.125 ;
        RECT 602.790 795.720 612.530 796.125 ;
        RECT 613.370 795.720 623.110 796.125 ;
        RECT 623.950 795.720 634.150 796.125 ;
        RECT 634.990 795.720 644.730 796.125 ;
        RECT 645.570 795.720 655.310 796.125 ;
        RECT 656.150 795.720 665.890 796.125 ;
        RECT 666.730 795.720 676.470 796.125 ;
        RECT 677.310 795.720 687.050 796.125 ;
        RECT 687.890 795.720 698.090 796.125 ;
        RECT 698.930 795.720 708.670 796.125 ;
        RECT 709.510 795.720 719.250 796.125 ;
        RECT 720.090 795.720 729.830 796.125 ;
        RECT 730.670 795.720 740.410 796.125 ;
        RECT 741.250 795.720 751.450 796.125 ;
        RECT 752.290 795.720 762.030 796.125 ;
        RECT 762.870 795.720 772.610 796.125 ;
        RECT 773.450 795.720 783.190 796.125 ;
        RECT 784.030 795.720 793.770 796.125 ;
        RECT 794.610 795.720 799.840 796.125 ;
        RECT 0.090 4.280 799.840 795.720 ;
        RECT 0.090 0.010 5.790 4.280 ;
        RECT 6.630 0.010 17.750 4.280 ;
        RECT 18.590 0.010 29.710 4.280 ;
        RECT 30.550 0.010 42.130 4.280 ;
        RECT 42.970 0.010 54.090 4.280 ;
        RECT 54.930 0.010 66.050 4.280 ;
        RECT 66.890 0.010 78.470 4.280 ;
        RECT 79.310 0.010 90.430 4.280 ;
        RECT 91.270 0.010 102.390 4.280 ;
        RECT 103.230 0.010 114.810 4.280 ;
        RECT 115.650 0.010 126.770 4.280 ;
        RECT 127.610 0.010 138.730 4.280 ;
        RECT 139.570 0.010 151.150 4.280 ;
        RECT 151.990 0.010 163.110 4.280 ;
        RECT 163.950 0.010 175.070 4.280 ;
        RECT 175.910 0.010 187.490 4.280 ;
        RECT 188.330 0.010 199.450 4.280 ;
        RECT 200.290 0.010 211.410 4.280 ;
        RECT 212.250 0.010 223.830 4.280 ;
        RECT 224.670 0.010 235.790 4.280 ;
        RECT 236.630 0.010 247.750 4.280 ;
        RECT 248.590 0.010 260.170 4.280 ;
        RECT 261.010 0.010 272.130 4.280 ;
        RECT 272.970 0.010 284.550 4.280 ;
        RECT 285.390 0.010 296.510 4.280 ;
        RECT 297.350 0.010 308.470 4.280 ;
        RECT 309.310 0.010 320.890 4.280 ;
        RECT 321.730 0.010 332.850 4.280 ;
        RECT 333.690 0.010 344.810 4.280 ;
        RECT 345.650 0.010 357.230 4.280 ;
        RECT 358.070 0.010 369.190 4.280 ;
        RECT 370.030 0.010 381.150 4.280 ;
        RECT 381.990 0.010 393.570 4.280 ;
        RECT 394.410 0.010 405.530 4.280 ;
        RECT 406.370 0.010 417.490 4.280 ;
        RECT 418.330 0.010 429.910 4.280 ;
        RECT 430.750 0.010 441.870 4.280 ;
        RECT 442.710 0.010 453.830 4.280 ;
        RECT 454.670 0.010 466.250 4.280 ;
        RECT 467.090 0.010 478.210 4.280 ;
        RECT 479.050 0.010 490.170 4.280 ;
        RECT 491.010 0.010 502.590 4.280 ;
        RECT 503.430 0.010 514.550 4.280 ;
        RECT 515.390 0.010 526.510 4.280 ;
        RECT 527.350 0.010 538.930 4.280 ;
        RECT 539.770 0.010 550.890 4.280 ;
        RECT 551.730 0.010 563.310 4.280 ;
        RECT 564.150 0.010 575.270 4.280 ;
        RECT 576.110 0.010 587.230 4.280 ;
        RECT 588.070 0.010 599.650 4.280 ;
        RECT 600.490 0.010 611.610 4.280 ;
        RECT 612.450 0.010 623.570 4.280 ;
        RECT 624.410 0.010 635.990 4.280 ;
        RECT 636.830 0.010 647.950 4.280 ;
        RECT 648.790 0.010 659.910 4.280 ;
        RECT 660.750 0.010 672.330 4.280 ;
        RECT 673.170 0.010 684.290 4.280 ;
        RECT 685.130 0.010 696.250 4.280 ;
        RECT 697.090 0.010 708.670 4.280 ;
        RECT 709.510 0.010 720.630 4.280 ;
        RECT 721.470 0.010 732.590 4.280 ;
        RECT 733.430 0.010 745.010 4.280 ;
        RECT 745.850 0.010 756.970 4.280 ;
        RECT 757.810 0.010 768.930 4.280 ;
        RECT 769.770 0.010 781.350 4.280 ;
        RECT 782.190 0.010 793.310 4.280 ;
        RECT 794.150 0.010 799.840 4.280 ;
      LAYER met3 ;
        RECT 0.065 795.240 795.600 796.105 ;
        RECT 0.065 793.920 796.000 795.240 ;
        RECT 4.400 792.520 796.000 793.920 ;
        RECT 0.065 789.840 796.000 792.520 ;
        RECT 0.065 788.440 795.600 789.840 ;
        RECT 0.065 783.040 796.000 788.440 ;
        RECT 0.065 781.680 795.600 783.040 ;
        RECT 4.400 781.640 795.600 781.680 ;
        RECT 4.400 780.280 796.000 781.640 ;
        RECT 0.065 776.240 796.000 780.280 ;
        RECT 0.065 774.840 795.600 776.240 ;
        RECT 0.065 768.760 796.000 774.840 ;
        RECT 4.400 767.360 795.600 768.760 ;
        RECT 0.065 761.960 796.000 767.360 ;
        RECT 0.065 760.560 795.600 761.960 ;
        RECT 0.065 756.520 796.000 760.560 ;
        RECT 4.400 755.160 796.000 756.520 ;
        RECT 4.400 755.120 795.600 755.160 ;
        RECT 0.065 753.760 795.600 755.120 ;
        RECT 0.065 748.360 796.000 753.760 ;
        RECT 0.065 746.960 795.600 748.360 ;
        RECT 0.065 744.280 796.000 746.960 ;
        RECT 4.400 742.880 796.000 744.280 ;
        RECT 0.065 740.880 796.000 742.880 ;
        RECT 0.065 739.480 795.600 740.880 ;
        RECT 0.065 734.080 796.000 739.480 ;
        RECT 0.065 732.680 795.600 734.080 ;
        RECT 0.065 731.360 796.000 732.680 ;
        RECT 4.400 729.960 796.000 731.360 ;
        RECT 0.065 727.280 796.000 729.960 ;
        RECT 0.065 725.880 795.600 727.280 ;
        RECT 0.065 720.480 796.000 725.880 ;
        RECT 0.065 719.120 795.600 720.480 ;
        RECT 4.400 719.080 795.600 719.120 ;
        RECT 4.400 717.720 796.000 719.080 ;
        RECT 0.065 713.680 796.000 717.720 ;
        RECT 0.065 712.280 795.600 713.680 ;
        RECT 0.065 706.880 796.000 712.280 ;
        RECT 4.400 706.200 796.000 706.880 ;
        RECT 4.400 705.480 795.600 706.200 ;
        RECT 0.065 704.800 795.600 705.480 ;
        RECT 0.065 699.400 796.000 704.800 ;
        RECT 0.065 698.000 795.600 699.400 ;
        RECT 0.065 693.960 796.000 698.000 ;
        RECT 4.400 692.600 796.000 693.960 ;
        RECT 4.400 692.560 795.600 692.600 ;
        RECT 0.065 691.200 795.600 692.560 ;
        RECT 0.065 685.800 796.000 691.200 ;
        RECT 0.065 684.400 795.600 685.800 ;
        RECT 0.065 681.720 796.000 684.400 ;
        RECT 4.400 680.320 796.000 681.720 ;
        RECT 0.065 678.320 796.000 680.320 ;
        RECT 0.065 676.920 795.600 678.320 ;
        RECT 0.065 671.520 796.000 676.920 ;
        RECT 0.065 670.120 795.600 671.520 ;
        RECT 0.065 668.800 796.000 670.120 ;
        RECT 4.400 667.400 796.000 668.800 ;
        RECT 0.065 664.720 796.000 667.400 ;
        RECT 0.065 663.320 795.600 664.720 ;
        RECT 0.065 657.920 796.000 663.320 ;
        RECT 0.065 656.560 795.600 657.920 ;
        RECT 4.400 656.520 795.600 656.560 ;
        RECT 4.400 655.160 796.000 656.520 ;
        RECT 0.065 651.120 796.000 655.160 ;
        RECT 0.065 649.720 795.600 651.120 ;
        RECT 0.065 644.320 796.000 649.720 ;
        RECT 4.400 643.640 796.000 644.320 ;
        RECT 4.400 642.920 795.600 643.640 ;
        RECT 0.065 642.240 795.600 642.920 ;
        RECT 0.065 636.840 796.000 642.240 ;
        RECT 0.065 635.440 795.600 636.840 ;
        RECT 0.065 631.400 796.000 635.440 ;
        RECT 4.400 630.040 796.000 631.400 ;
        RECT 4.400 630.000 795.600 630.040 ;
        RECT 0.065 628.640 795.600 630.000 ;
        RECT 0.065 623.240 796.000 628.640 ;
        RECT 0.065 621.840 795.600 623.240 ;
        RECT 0.065 619.160 796.000 621.840 ;
        RECT 4.400 617.760 796.000 619.160 ;
        RECT 0.065 615.760 796.000 617.760 ;
        RECT 0.065 614.360 795.600 615.760 ;
        RECT 0.065 608.960 796.000 614.360 ;
        RECT 0.065 607.560 795.600 608.960 ;
        RECT 0.065 606.920 796.000 607.560 ;
        RECT 4.400 605.520 796.000 606.920 ;
        RECT 0.065 602.160 796.000 605.520 ;
        RECT 0.065 600.760 795.600 602.160 ;
        RECT 0.065 595.360 796.000 600.760 ;
        RECT 0.065 594.000 795.600 595.360 ;
        RECT 4.400 593.960 795.600 594.000 ;
        RECT 4.400 592.600 796.000 593.960 ;
        RECT 0.065 587.880 796.000 592.600 ;
        RECT 0.065 586.480 795.600 587.880 ;
        RECT 0.065 581.760 796.000 586.480 ;
        RECT 4.400 581.080 796.000 581.760 ;
        RECT 4.400 580.360 795.600 581.080 ;
        RECT 0.065 579.680 795.600 580.360 ;
        RECT 0.065 574.280 796.000 579.680 ;
        RECT 0.065 572.880 795.600 574.280 ;
        RECT 0.065 568.840 796.000 572.880 ;
        RECT 4.400 567.480 796.000 568.840 ;
        RECT 4.400 567.440 795.600 567.480 ;
        RECT 0.065 566.080 795.600 567.440 ;
        RECT 0.065 560.680 796.000 566.080 ;
        RECT 0.065 559.280 795.600 560.680 ;
        RECT 0.065 556.600 796.000 559.280 ;
        RECT 4.400 555.200 796.000 556.600 ;
        RECT 0.065 553.200 796.000 555.200 ;
        RECT 0.065 551.800 795.600 553.200 ;
        RECT 0.065 546.400 796.000 551.800 ;
        RECT 0.065 545.000 795.600 546.400 ;
        RECT 0.065 544.360 796.000 545.000 ;
        RECT 4.400 542.960 796.000 544.360 ;
        RECT 0.065 539.600 796.000 542.960 ;
        RECT 0.065 538.200 795.600 539.600 ;
        RECT 0.065 532.800 796.000 538.200 ;
        RECT 0.065 531.440 795.600 532.800 ;
        RECT 4.400 531.400 795.600 531.440 ;
        RECT 4.400 530.040 796.000 531.400 ;
        RECT 0.065 525.320 796.000 530.040 ;
        RECT 0.065 523.920 795.600 525.320 ;
        RECT 0.065 519.200 796.000 523.920 ;
        RECT 4.400 518.520 796.000 519.200 ;
        RECT 4.400 517.800 795.600 518.520 ;
        RECT 0.065 517.120 795.600 517.800 ;
        RECT 0.065 511.720 796.000 517.120 ;
        RECT 0.065 510.320 795.600 511.720 ;
        RECT 0.065 506.960 796.000 510.320 ;
        RECT 4.400 505.560 796.000 506.960 ;
        RECT 0.065 504.920 796.000 505.560 ;
        RECT 0.065 503.520 795.600 504.920 ;
        RECT 0.065 498.120 796.000 503.520 ;
        RECT 0.065 496.720 795.600 498.120 ;
        RECT 0.065 494.040 796.000 496.720 ;
        RECT 4.400 492.640 796.000 494.040 ;
        RECT 0.065 490.640 796.000 492.640 ;
        RECT 0.065 489.240 795.600 490.640 ;
        RECT 0.065 483.840 796.000 489.240 ;
        RECT 0.065 482.440 795.600 483.840 ;
        RECT 0.065 481.800 796.000 482.440 ;
        RECT 4.400 480.400 796.000 481.800 ;
        RECT 0.065 477.040 796.000 480.400 ;
        RECT 0.065 475.640 795.600 477.040 ;
        RECT 0.065 470.240 796.000 475.640 ;
        RECT 0.065 468.880 795.600 470.240 ;
        RECT 4.400 468.840 795.600 468.880 ;
        RECT 4.400 467.480 796.000 468.840 ;
        RECT 0.065 462.760 796.000 467.480 ;
        RECT 0.065 461.360 795.600 462.760 ;
        RECT 0.065 456.640 796.000 461.360 ;
        RECT 4.400 455.960 796.000 456.640 ;
        RECT 4.400 455.240 795.600 455.960 ;
        RECT 0.065 454.560 795.600 455.240 ;
        RECT 0.065 449.160 796.000 454.560 ;
        RECT 0.065 447.760 795.600 449.160 ;
        RECT 0.065 444.400 796.000 447.760 ;
        RECT 4.400 443.000 796.000 444.400 ;
        RECT 0.065 442.360 796.000 443.000 ;
        RECT 0.065 440.960 795.600 442.360 ;
        RECT 0.065 435.560 796.000 440.960 ;
        RECT 0.065 434.160 795.600 435.560 ;
        RECT 0.065 431.480 796.000 434.160 ;
        RECT 4.400 430.080 796.000 431.480 ;
        RECT 0.065 428.080 796.000 430.080 ;
        RECT 0.065 426.680 795.600 428.080 ;
        RECT 0.065 421.280 796.000 426.680 ;
        RECT 0.065 419.880 795.600 421.280 ;
        RECT 0.065 419.240 796.000 419.880 ;
        RECT 4.400 417.840 796.000 419.240 ;
        RECT 0.065 414.480 796.000 417.840 ;
        RECT 0.065 413.080 795.600 414.480 ;
        RECT 0.065 407.680 796.000 413.080 ;
        RECT 0.065 407.000 795.600 407.680 ;
        RECT 4.400 406.280 795.600 407.000 ;
        RECT 4.400 405.600 796.000 406.280 ;
        RECT 0.065 400.200 796.000 405.600 ;
        RECT 0.065 398.800 795.600 400.200 ;
        RECT 0.065 394.080 796.000 398.800 ;
        RECT 4.400 393.400 796.000 394.080 ;
        RECT 4.400 392.680 795.600 393.400 ;
        RECT 0.065 392.000 795.600 392.680 ;
        RECT 0.065 386.600 796.000 392.000 ;
        RECT 0.065 385.200 795.600 386.600 ;
        RECT 0.065 381.840 796.000 385.200 ;
        RECT 4.400 380.440 796.000 381.840 ;
        RECT 0.065 379.800 796.000 380.440 ;
        RECT 0.065 378.400 795.600 379.800 ;
        RECT 0.065 372.320 796.000 378.400 ;
        RECT 0.065 370.920 795.600 372.320 ;
        RECT 0.065 368.920 796.000 370.920 ;
        RECT 4.400 367.520 796.000 368.920 ;
        RECT 0.065 365.520 796.000 367.520 ;
        RECT 0.065 364.120 795.600 365.520 ;
        RECT 0.065 358.720 796.000 364.120 ;
        RECT 0.065 357.320 795.600 358.720 ;
        RECT 0.065 356.680 796.000 357.320 ;
        RECT 4.400 355.280 796.000 356.680 ;
        RECT 0.065 351.920 796.000 355.280 ;
        RECT 0.065 350.520 795.600 351.920 ;
        RECT 0.065 345.120 796.000 350.520 ;
        RECT 0.065 344.440 795.600 345.120 ;
        RECT 4.400 343.720 795.600 344.440 ;
        RECT 4.400 343.040 796.000 343.720 ;
        RECT 0.065 337.640 796.000 343.040 ;
        RECT 0.065 336.240 795.600 337.640 ;
        RECT 0.065 331.520 796.000 336.240 ;
        RECT 4.400 330.840 796.000 331.520 ;
        RECT 4.400 330.120 795.600 330.840 ;
        RECT 0.065 329.440 795.600 330.120 ;
        RECT 0.065 324.040 796.000 329.440 ;
        RECT 0.065 322.640 795.600 324.040 ;
        RECT 0.065 319.280 796.000 322.640 ;
        RECT 4.400 317.880 796.000 319.280 ;
        RECT 0.065 317.240 796.000 317.880 ;
        RECT 0.065 315.840 795.600 317.240 ;
        RECT 0.065 309.760 796.000 315.840 ;
        RECT 0.065 308.360 795.600 309.760 ;
        RECT 0.065 307.040 796.000 308.360 ;
        RECT 4.400 305.640 796.000 307.040 ;
        RECT 0.065 302.960 796.000 305.640 ;
        RECT 0.065 301.560 795.600 302.960 ;
        RECT 0.065 296.160 796.000 301.560 ;
        RECT 0.065 294.760 795.600 296.160 ;
        RECT 0.065 294.120 796.000 294.760 ;
        RECT 4.400 292.720 796.000 294.120 ;
        RECT 0.065 289.360 796.000 292.720 ;
        RECT 0.065 287.960 795.600 289.360 ;
        RECT 0.065 282.560 796.000 287.960 ;
        RECT 0.065 281.880 795.600 282.560 ;
        RECT 4.400 281.160 795.600 281.880 ;
        RECT 4.400 280.480 796.000 281.160 ;
        RECT 0.065 275.080 796.000 280.480 ;
        RECT 0.065 273.680 795.600 275.080 ;
        RECT 0.065 268.960 796.000 273.680 ;
        RECT 4.400 268.280 796.000 268.960 ;
        RECT 4.400 267.560 795.600 268.280 ;
        RECT 0.065 266.880 795.600 267.560 ;
        RECT 0.065 261.480 796.000 266.880 ;
        RECT 0.065 260.080 795.600 261.480 ;
        RECT 0.065 256.720 796.000 260.080 ;
        RECT 4.400 255.320 796.000 256.720 ;
        RECT 0.065 254.680 796.000 255.320 ;
        RECT 0.065 253.280 795.600 254.680 ;
        RECT 0.065 247.200 796.000 253.280 ;
        RECT 0.065 245.800 795.600 247.200 ;
        RECT 0.065 244.480 796.000 245.800 ;
        RECT 4.400 243.080 796.000 244.480 ;
        RECT 0.065 240.400 796.000 243.080 ;
        RECT 0.065 239.000 795.600 240.400 ;
        RECT 0.065 233.600 796.000 239.000 ;
        RECT 0.065 232.200 795.600 233.600 ;
        RECT 0.065 231.560 796.000 232.200 ;
        RECT 4.400 230.160 796.000 231.560 ;
        RECT 0.065 226.800 796.000 230.160 ;
        RECT 0.065 225.400 795.600 226.800 ;
        RECT 0.065 220.000 796.000 225.400 ;
        RECT 0.065 219.320 795.600 220.000 ;
        RECT 4.400 218.600 795.600 219.320 ;
        RECT 4.400 217.920 796.000 218.600 ;
        RECT 0.065 212.520 796.000 217.920 ;
        RECT 0.065 211.120 795.600 212.520 ;
        RECT 0.065 207.080 796.000 211.120 ;
        RECT 4.400 205.720 796.000 207.080 ;
        RECT 4.400 205.680 795.600 205.720 ;
        RECT 0.065 204.320 795.600 205.680 ;
        RECT 0.065 198.920 796.000 204.320 ;
        RECT 0.065 197.520 795.600 198.920 ;
        RECT 0.065 194.160 796.000 197.520 ;
        RECT 4.400 192.760 796.000 194.160 ;
        RECT 0.065 192.120 796.000 192.760 ;
        RECT 0.065 190.720 795.600 192.120 ;
        RECT 0.065 184.640 796.000 190.720 ;
        RECT 0.065 183.240 795.600 184.640 ;
        RECT 0.065 181.920 796.000 183.240 ;
        RECT 4.400 180.520 796.000 181.920 ;
        RECT 0.065 177.840 796.000 180.520 ;
        RECT 0.065 176.440 795.600 177.840 ;
        RECT 0.065 171.040 796.000 176.440 ;
        RECT 0.065 169.640 795.600 171.040 ;
        RECT 0.065 169.000 796.000 169.640 ;
        RECT 4.400 167.600 796.000 169.000 ;
        RECT 0.065 164.240 796.000 167.600 ;
        RECT 0.065 162.840 795.600 164.240 ;
        RECT 0.065 156.760 796.000 162.840 ;
        RECT 4.400 155.360 795.600 156.760 ;
        RECT 0.065 149.960 796.000 155.360 ;
        RECT 0.065 148.560 795.600 149.960 ;
        RECT 0.065 144.520 796.000 148.560 ;
        RECT 4.400 143.160 796.000 144.520 ;
        RECT 4.400 143.120 795.600 143.160 ;
        RECT 0.065 141.760 795.600 143.120 ;
        RECT 0.065 136.360 796.000 141.760 ;
        RECT 0.065 134.960 795.600 136.360 ;
        RECT 0.065 131.600 796.000 134.960 ;
        RECT 4.400 130.200 796.000 131.600 ;
        RECT 0.065 129.560 796.000 130.200 ;
        RECT 0.065 128.160 795.600 129.560 ;
        RECT 0.065 122.080 796.000 128.160 ;
        RECT 0.065 120.680 795.600 122.080 ;
        RECT 0.065 119.360 796.000 120.680 ;
        RECT 4.400 117.960 796.000 119.360 ;
        RECT 0.065 115.280 796.000 117.960 ;
        RECT 0.065 113.880 795.600 115.280 ;
        RECT 0.065 108.480 796.000 113.880 ;
        RECT 0.065 107.120 795.600 108.480 ;
        RECT 4.400 107.080 795.600 107.120 ;
        RECT 4.400 105.720 796.000 107.080 ;
        RECT 0.065 101.680 796.000 105.720 ;
        RECT 0.065 100.280 795.600 101.680 ;
        RECT 0.065 94.200 796.000 100.280 ;
        RECT 4.400 92.800 795.600 94.200 ;
        RECT 0.065 87.400 796.000 92.800 ;
        RECT 0.065 86.000 795.600 87.400 ;
        RECT 0.065 81.960 796.000 86.000 ;
        RECT 4.400 80.600 796.000 81.960 ;
        RECT 4.400 80.560 795.600 80.600 ;
        RECT 0.065 79.200 795.600 80.560 ;
        RECT 0.065 73.800 796.000 79.200 ;
        RECT 0.065 72.400 795.600 73.800 ;
        RECT 0.065 69.040 796.000 72.400 ;
        RECT 4.400 67.640 796.000 69.040 ;
        RECT 0.065 67.000 796.000 67.640 ;
        RECT 0.065 65.600 795.600 67.000 ;
        RECT 0.065 59.520 796.000 65.600 ;
        RECT 0.065 58.120 795.600 59.520 ;
        RECT 0.065 56.800 796.000 58.120 ;
        RECT 4.400 55.400 796.000 56.800 ;
        RECT 0.065 52.720 796.000 55.400 ;
        RECT 0.065 51.320 795.600 52.720 ;
        RECT 0.065 45.920 796.000 51.320 ;
        RECT 0.065 44.560 795.600 45.920 ;
        RECT 4.400 44.520 795.600 44.560 ;
        RECT 4.400 43.160 796.000 44.520 ;
        RECT 0.065 39.120 796.000 43.160 ;
        RECT 0.065 37.720 795.600 39.120 ;
        RECT 0.065 31.640 796.000 37.720 ;
        RECT 4.400 30.240 795.600 31.640 ;
        RECT 0.065 24.840 796.000 30.240 ;
        RECT 0.065 23.440 795.600 24.840 ;
        RECT 0.065 19.400 796.000 23.440 ;
        RECT 4.400 18.040 796.000 19.400 ;
        RECT 4.400 18.000 795.600 18.040 ;
        RECT 0.065 16.640 795.600 18.000 ;
        RECT 0.065 11.240 796.000 16.640 ;
        RECT 0.065 9.840 795.600 11.240 ;
        RECT 0.065 7.160 796.000 9.840 ;
        RECT 4.400 5.760 796.000 7.160 ;
        RECT 0.065 4.440 796.000 5.760 ;
        RECT 0.065 3.040 795.600 4.440 ;
        RECT 0.065 0.175 796.000 3.040 ;
      LAYER met4 ;
        RECT 0.295 10.240 20.640 784.545 ;
        RECT 23.040 10.480 23.940 784.545 ;
        RECT 26.340 10.480 27.240 784.545 ;
        RECT 29.640 10.480 30.540 784.545 ;
        RECT 32.940 10.480 97.440 784.545 ;
        RECT 23.040 10.240 97.440 10.480 ;
        RECT 99.840 10.480 100.740 784.545 ;
        RECT 103.140 10.480 104.040 784.545 ;
        RECT 106.440 10.480 107.340 784.545 ;
        RECT 109.740 10.480 174.240 784.545 ;
        RECT 99.840 10.240 174.240 10.480 ;
        RECT 176.640 10.480 177.540 784.545 ;
        RECT 179.940 10.480 180.840 784.545 ;
        RECT 183.240 10.480 184.140 784.545 ;
        RECT 186.540 10.480 251.040 784.545 ;
        RECT 176.640 10.240 251.040 10.480 ;
        RECT 253.440 10.480 254.340 784.545 ;
        RECT 256.740 10.480 257.640 784.545 ;
        RECT 260.040 10.480 260.940 784.545 ;
        RECT 263.340 10.480 327.840 784.545 ;
        RECT 253.440 10.240 327.840 10.480 ;
        RECT 330.240 10.480 331.140 784.545 ;
        RECT 333.540 10.480 334.440 784.545 ;
        RECT 336.840 10.480 337.740 784.545 ;
        RECT 340.140 10.480 404.640 784.545 ;
        RECT 330.240 10.240 404.640 10.480 ;
        RECT 407.040 10.480 407.940 784.545 ;
        RECT 410.340 10.480 411.240 784.545 ;
        RECT 413.640 10.480 414.540 784.545 ;
        RECT 416.940 10.480 481.440 784.545 ;
        RECT 407.040 10.240 481.440 10.480 ;
        RECT 483.840 10.480 484.740 784.545 ;
        RECT 487.140 10.480 488.040 784.545 ;
        RECT 490.440 10.480 491.340 784.545 ;
        RECT 493.740 10.480 558.240 784.545 ;
        RECT 483.840 10.240 558.240 10.480 ;
        RECT 560.640 10.480 561.540 784.545 ;
        RECT 563.940 10.480 564.840 784.545 ;
        RECT 567.240 10.480 568.140 784.545 ;
        RECT 570.540 10.480 635.040 784.545 ;
        RECT 560.640 10.240 635.040 10.480 ;
        RECT 637.440 10.480 638.340 784.545 ;
        RECT 640.740 10.480 641.640 784.545 ;
        RECT 644.040 10.480 644.940 784.545 ;
        RECT 647.340 10.480 711.840 784.545 ;
        RECT 637.440 10.240 711.840 10.480 ;
        RECT 714.240 10.480 715.140 784.545 ;
        RECT 717.540 10.480 718.440 784.545 ;
        RECT 720.840 10.480 721.740 784.545 ;
        RECT 724.140 10.480 785.385 784.545 ;
        RECT 714.240 10.240 785.385 10.480 ;
        RECT 0.295 0.175 785.385 10.240 ;
  END
END wrapper_sha1
END LIBRARY

