VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapper_sha1
  CLASS BLOCK ;
  FOREIGN wrapper_sha1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 673.055 BY 683.775 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 679.775 58.330 683.775 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 2.760 673.055 3.360 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 180.920 673.055 181.520 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 198.600 673.055 199.200 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 216.280 673.055 216.880 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 234.640 673.055 235.240 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 252.320 673.055 252.920 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 270.000 673.055 270.600 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 287.680 673.055 288.280 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 306.040 673.055 306.640 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 323.720 673.055 324.320 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 341.400 673.055 342.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 20.440 673.055 21.040 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 359.080 673.055 359.680 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 377.440 673.055 378.040 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 395.120 673.055 395.720 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 412.800 673.055 413.400 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 430.480 673.055 431.080 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 448.840 673.055 449.440 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 466.520 673.055 467.120 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 484.200 673.055 484.800 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 501.880 673.055 502.480 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 520.240 673.055 520.840 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 38.120 673.055 38.720 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 537.920 673.055 538.520 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 555.600 673.055 556.200 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 573.280 673.055 573.880 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 591.640 673.055 592.240 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 609.320 673.055 609.920 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 627.000 673.055 627.600 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 644.680 673.055 645.280 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 663.040 673.055 663.640 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 55.800 673.055 56.400 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 73.480 673.055 74.080 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 91.840 673.055 92.440 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 109.520 673.055 110.120 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 127.200 673.055 127.800 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 144.880 673.055 145.480 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 163.240 673.055 163.840 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 14.320 673.055 14.920 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 192.480 673.055 193.080 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 210.840 673.055 211.440 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 228.520 673.055 229.120 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 246.200 673.055 246.800 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 263.880 673.055 264.480 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 282.240 673.055 282.840 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 299.920 673.055 300.520 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 317.600 673.055 318.200 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 335.280 673.055 335.880 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 353.640 673.055 354.240 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 32.000 673.055 32.600 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 371.320 673.055 371.920 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 389.000 673.055 389.600 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 406.680 673.055 407.280 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 425.040 673.055 425.640 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 442.720 673.055 443.320 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 460.400 673.055 461.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 478.080 673.055 478.680 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 496.440 673.055 497.040 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 514.120 673.055 514.720 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 531.800 673.055 532.400 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 49.680 673.055 50.280 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 549.480 673.055 550.080 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 567.840 673.055 568.440 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 585.520 673.055 586.120 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 603.200 673.055 603.800 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 620.880 673.055 621.480 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 639.240 673.055 639.840 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 656.920 673.055 657.520 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 674.600 673.055 675.200 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 68.040 673.055 68.640 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 85.720 673.055 86.320 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 103.400 673.055 104.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 121.080 673.055 121.680 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 139.440 673.055 140.040 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 157.120 673.055 157.720 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 174.800 673.055 175.400 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 8.200 673.055 8.800 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 187.040 673.055 187.640 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 204.720 673.055 205.320 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 222.400 673.055 223.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 240.080 673.055 240.680 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 258.440 673.055 259.040 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 276.120 673.055 276.720 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 293.800 673.055 294.400 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 311.480 673.055 312.080 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 329.840 673.055 330.440 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 347.520 673.055 348.120 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 25.880 673.055 26.480 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 365.200 673.055 365.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 382.880 673.055 383.480 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 401.240 673.055 401.840 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 418.920 673.055 419.520 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 436.600 673.055 437.200 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 454.280 673.055 454.880 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 472.640 673.055 473.240 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 490.320 673.055 490.920 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 508.000 673.055 508.600 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 525.680 673.055 526.280 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 44.240 673.055 44.840 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 544.040 673.055 544.640 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 561.720 673.055 562.320 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 579.400 673.055 580.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 597.080 673.055 597.680 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 615.440 673.055 616.040 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 633.120 673.055 633.720 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 650.800 673.055 651.400 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 668.480 673.055 669.080 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 61.920 673.055 62.520 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 79.600 673.055 80.200 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 97.280 673.055 97.880 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 115.640 673.055 116.240 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 133.320 673.055 133.920 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 151.000 673.055 151.600 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 168.680 673.055 169.280 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 0.000 667.830 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.055 680.720 673.055 681.320 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.000 4.000 678.600 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 0.000 253.830 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 0.000 305.350 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 0.000 336.630 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 0.000 470.950 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 0.000 481.530 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 0.000 491.650 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 0.000 522.930 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 0.000 533.050 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 0.000 543.630 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 0.000 553.750 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 0.000 564.330 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 0.000 574.450 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 0.000 585.030 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 0.000 595.150 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 0.000 615.850 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 0.000 626.430 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 0.000 636.550 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.850 0.000 647.130 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 0.000 419.430 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.800 4.000 447.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.200 4.000 467.800 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.080 4.000 478.680 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 509.360 4.000 509.960 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 4.000 541.920 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.600 4.000 352.200 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 551.520 4.000 552.120 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 562.400 4.000 563.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.680 4.000 594.280 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 604.560 4.000 605.160 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.760 4.000 615.360 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.720 4.000 647.320 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 362.480 4.000 363.080 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.920 4.000 657.520 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.800 4.000 668.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.760 4.000 394.360 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.920 4.000 436.520 ;
    END
  END la_oenb[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 679.775 4.510 683.775 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 679.775 13.250 683.775 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 679.775 49.130 683.775 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 679.775 102.950 683.775 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 679.775 192.650 683.775 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 679.775 201.850 683.775 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 679.775 210.590 683.775 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 679.775 219.790 683.775 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 679.775 228.530 683.775 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 679.775 237.730 683.775 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 679.775 246.470 683.775 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 679.775 255.670 683.775 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 679.775 264.410 683.775 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 679.775 273.610 683.775 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 679.775 112.150 683.775 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 679.775 282.350 683.775 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 679.775 291.550 683.775 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 679.775 300.290 683.775 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 679.775 309.490 683.775 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 679.775 318.230 683.775 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 679.775 327.430 683.775 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 679.775 336.170 683.775 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 679.775 345.370 683.775 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 679.775 354.110 683.775 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 679.775 363.310 683.775 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 679.775 120.890 683.775 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 679.775 372.050 683.775 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 679.775 381.250 683.775 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 679.775 130.090 683.775 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 679.775 138.830 683.775 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 679.775 148.030 683.775 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 679.775 156.770 683.775 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 679.775 165.970 683.775 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 679.775 174.710 683.775 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 679.775 183.910 683.775 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 679.775 31.190 683.775 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 679.775 389.990 683.775 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 679.775 479.690 683.775 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 679.775 488.890 683.775 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 679.775 497.630 683.775 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 679.775 506.830 683.775 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 679.775 515.570 683.775 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 679.775 524.770 683.775 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 679.775 533.510 683.775 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 679.775 542.710 683.775 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 679.775 551.450 683.775 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 679.775 560.650 683.775 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 679.775 399.190 683.775 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 679.775 569.390 683.775 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 679.775 578.590 683.775 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 679.775 587.330 683.775 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 679.775 596.530 683.775 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 679.775 605.270 683.775 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 679.775 614.470 683.775 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 679.775 623.210 683.775 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 679.775 632.410 683.775 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 679.775 641.150 683.775 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 679.775 650.350 683.775 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 679.775 407.930 683.775 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 679.775 659.090 683.775 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.010 679.775 668.290 683.775 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 679.775 417.130 683.775 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 679.775 425.870 683.775 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 679.775 435.070 683.775 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 679.775 443.810 683.775 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 679.775 453.010 683.775 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 679.775 461.750 683.775 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 679.775 470.950 683.775 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.280 4.000 267.880 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 679.775 67.070 683.775 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 679.775 76.270 683.775 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 679.775 85.010 683.775 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 679.775 94.210 683.775 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 679.775 22.450 683.775 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 679.775 40.390 683.775 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 672.080 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 672.080 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 672.080 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 672.080 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 672.080 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 639.210 667.460 640.810 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 486.030 667.460 487.630 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 332.850 667.460 334.450 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 179.670 667.460 181.270 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 667.460 28.090 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 672.080 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 672.080 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 672.080 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 672.080 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 562.620 667.460 564.220 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 409.440 667.460 411.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 256.260 667.460 257.860 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 667.460 104.680 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.740 10.880 640.340 671.840 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 671.840 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 671.840 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 671.840 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 671.840 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 642.750 667.460 644.350 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 489.570 667.460 491.170 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 336.390 667.460 337.990 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 183.210 667.460 184.810 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 30.030 667.460 31.630 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.940 10.880 563.540 671.840 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 671.840 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 671.840 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 671.840 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 566.160 667.460 567.760 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 412.980 667.460 414.580 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 259.800 667.460 261.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 106.620 667.460 108.220 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 642.040 10.880 643.640 671.840 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 488.440 10.880 490.040 671.840 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 671.840 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 671.840 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 671.840 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 646.050 667.460 647.650 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 492.870 667.460 494.470 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 339.690 667.460 341.290 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 186.510 667.460 188.110 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 33.330 667.460 34.930 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 565.240 10.880 566.840 671.840 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.640 10.880 413.240 671.840 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 671.840 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 671.840 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 569.460 667.460 571.060 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 416.280 667.460 417.880 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 263.100 667.460 264.700 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 109.920 667.460 111.520 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 645.340 10.880 646.940 671.840 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 491.740 10.880 493.340 671.840 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 671.840 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 671.840 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 671.840 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 649.350 667.460 650.950 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 496.170 667.460 497.770 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 342.990 667.460 344.590 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 189.810 667.460 191.410 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 36.630 667.460 38.230 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 568.540 10.880 570.140 671.840 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 414.940 10.880 416.540 671.840 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 671.840 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 671.840 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 572.760 667.460 574.360 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 419.580 667.460 421.180 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 266.400 667.460 268.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 113.220 667.460 114.820 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 0.605 0.085 672.375 682.635 ;
      LAYER met1 ;
        RECT 0.070 0.040 672.910 683.700 ;
      LAYER met2 ;
        RECT 0.090 679.495 3.950 683.730 ;
        RECT 4.790 679.495 12.690 683.730 ;
        RECT 13.530 679.495 21.890 683.730 ;
        RECT 22.730 679.495 30.630 683.730 ;
        RECT 31.470 679.495 39.830 683.730 ;
        RECT 40.670 679.495 48.570 683.730 ;
        RECT 49.410 679.495 57.770 683.730 ;
        RECT 58.610 679.495 66.510 683.730 ;
        RECT 67.350 679.495 75.710 683.730 ;
        RECT 76.550 679.495 84.450 683.730 ;
        RECT 85.290 679.495 93.650 683.730 ;
        RECT 94.490 679.495 102.390 683.730 ;
        RECT 103.230 679.495 111.590 683.730 ;
        RECT 112.430 679.495 120.330 683.730 ;
        RECT 121.170 679.495 129.530 683.730 ;
        RECT 130.370 679.495 138.270 683.730 ;
        RECT 139.110 679.495 147.470 683.730 ;
        RECT 148.310 679.495 156.210 683.730 ;
        RECT 157.050 679.495 165.410 683.730 ;
        RECT 166.250 679.495 174.150 683.730 ;
        RECT 174.990 679.495 183.350 683.730 ;
        RECT 184.190 679.495 192.090 683.730 ;
        RECT 192.930 679.495 201.290 683.730 ;
        RECT 202.130 679.495 210.030 683.730 ;
        RECT 210.870 679.495 219.230 683.730 ;
        RECT 220.070 679.495 227.970 683.730 ;
        RECT 228.810 679.495 237.170 683.730 ;
        RECT 238.010 679.495 245.910 683.730 ;
        RECT 246.750 679.495 255.110 683.730 ;
        RECT 255.950 679.495 263.850 683.730 ;
        RECT 264.690 679.495 273.050 683.730 ;
        RECT 273.890 679.495 281.790 683.730 ;
        RECT 282.630 679.495 290.990 683.730 ;
        RECT 291.830 679.495 299.730 683.730 ;
        RECT 300.570 679.495 308.930 683.730 ;
        RECT 309.770 679.495 317.670 683.730 ;
        RECT 318.510 679.495 326.870 683.730 ;
        RECT 327.710 679.495 335.610 683.730 ;
        RECT 336.450 679.495 344.810 683.730 ;
        RECT 345.650 679.495 353.550 683.730 ;
        RECT 354.390 679.495 362.750 683.730 ;
        RECT 363.590 679.495 371.490 683.730 ;
        RECT 372.330 679.495 380.690 683.730 ;
        RECT 381.530 679.495 389.430 683.730 ;
        RECT 390.270 679.495 398.630 683.730 ;
        RECT 399.470 679.495 407.370 683.730 ;
        RECT 408.210 679.495 416.570 683.730 ;
        RECT 417.410 679.495 425.310 683.730 ;
        RECT 426.150 679.495 434.510 683.730 ;
        RECT 435.350 679.495 443.250 683.730 ;
        RECT 444.090 679.495 452.450 683.730 ;
        RECT 453.290 679.495 461.190 683.730 ;
        RECT 462.030 679.495 470.390 683.730 ;
        RECT 471.230 679.495 479.130 683.730 ;
        RECT 479.970 679.495 488.330 683.730 ;
        RECT 489.170 679.495 497.070 683.730 ;
        RECT 497.910 679.495 506.270 683.730 ;
        RECT 507.110 679.495 515.010 683.730 ;
        RECT 515.850 679.495 524.210 683.730 ;
        RECT 525.050 679.495 532.950 683.730 ;
        RECT 533.790 679.495 542.150 683.730 ;
        RECT 542.990 679.495 550.890 683.730 ;
        RECT 551.730 679.495 560.090 683.730 ;
        RECT 560.930 679.495 568.830 683.730 ;
        RECT 569.670 679.495 578.030 683.730 ;
        RECT 578.870 679.495 586.770 683.730 ;
        RECT 587.610 679.495 595.970 683.730 ;
        RECT 596.810 679.495 604.710 683.730 ;
        RECT 605.550 679.495 613.910 683.730 ;
        RECT 614.750 679.495 622.650 683.730 ;
        RECT 623.490 679.495 631.850 683.730 ;
        RECT 632.690 679.495 640.590 683.730 ;
        RECT 641.430 679.495 649.790 683.730 ;
        RECT 650.630 679.495 658.530 683.730 ;
        RECT 659.370 679.495 667.730 683.730 ;
        RECT 668.570 679.495 672.890 683.730 ;
        RECT 0.090 4.280 672.890 679.495 ;
        RECT 0.090 0.010 4.870 4.280 ;
        RECT 5.710 0.010 14.990 4.280 ;
        RECT 15.830 0.010 25.570 4.280 ;
        RECT 26.410 0.010 35.690 4.280 ;
        RECT 36.530 0.010 46.270 4.280 ;
        RECT 47.110 0.010 56.390 4.280 ;
        RECT 57.230 0.010 66.970 4.280 ;
        RECT 67.810 0.010 77.090 4.280 ;
        RECT 77.930 0.010 87.670 4.280 ;
        RECT 88.510 0.010 97.790 4.280 ;
        RECT 98.630 0.010 108.370 4.280 ;
        RECT 109.210 0.010 118.490 4.280 ;
        RECT 119.330 0.010 129.070 4.280 ;
        RECT 129.910 0.010 139.190 4.280 ;
        RECT 140.030 0.010 149.770 4.280 ;
        RECT 150.610 0.010 159.890 4.280 ;
        RECT 160.730 0.010 170.470 4.280 ;
        RECT 171.310 0.010 180.590 4.280 ;
        RECT 181.430 0.010 191.170 4.280 ;
        RECT 192.010 0.010 201.290 4.280 ;
        RECT 202.130 0.010 211.870 4.280 ;
        RECT 212.710 0.010 221.990 4.280 ;
        RECT 222.830 0.010 232.570 4.280 ;
        RECT 233.410 0.010 242.690 4.280 ;
        RECT 243.530 0.010 253.270 4.280 ;
        RECT 254.110 0.010 263.390 4.280 ;
        RECT 264.230 0.010 273.970 4.280 ;
        RECT 274.810 0.010 284.090 4.280 ;
        RECT 284.930 0.010 294.670 4.280 ;
        RECT 295.510 0.010 304.790 4.280 ;
        RECT 305.630 0.010 315.370 4.280 ;
        RECT 316.210 0.010 325.490 4.280 ;
        RECT 326.330 0.010 336.070 4.280 ;
        RECT 336.910 0.010 346.190 4.280 ;
        RECT 347.030 0.010 356.770 4.280 ;
        RECT 357.610 0.010 366.890 4.280 ;
        RECT 367.730 0.010 377.470 4.280 ;
        RECT 378.310 0.010 387.590 4.280 ;
        RECT 388.430 0.010 398.170 4.280 ;
        RECT 399.010 0.010 408.290 4.280 ;
        RECT 409.130 0.010 418.870 4.280 ;
        RECT 419.710 0.010 428.990 4.280 ;
        RECT 429.830 0.010 439.570 4.280 ;
        RECT 440.410 0.010 449.690 4.280 ;
        RECT 450.530 0.010 460.270 4.280 ;
        RECT 461.110 0.010 470.390 4.280 ;
        RECT 471.230 0.010 480.970 4.280 ;
        RECT 481.810 0.010 491.090 4.280 ;
        RECT 491.930 0.010 501.670 4.280 ;
        RECT 502.510 0.010 511.790 4.280 ;
        RECT 512.630 0.010 522.370 4.280 ;
        RECT 523.210 0.010 532.490 4.280 ;
        RECT 533.330 0.010 543.070 4.280 ;
        RECT 543.910 0.010 553.190 4.280 ;
        RECT 554.030 0.010 563.770 4.280 ;
        RECT 564.610 0.010 573.890 4.280 ;
        RECT 574.730 0.010 584.470 4.280 ;
        RECT 585.310 0.010 594.590 4.280 ;
        RECT 595.430 0.010 605.170 4.280 ;
        RECT 606.010 0.010 615.290 4.280 ;
        RECT 616.130 0.010 625.870 4.280 ;
        RECT 626.710 0.010 635.990 4.280 ;
        RECT 636.830 0.010 646.570 4.280 ;
        RECT 647.410 0.010 656.690 4.280 ;
        RECT 657.530 0.010 667.270 4.280 ;
        RECT 668.110 0.010 672.890 4.280 ;
      LAYER met3 ;
        RECT 0.065 680.320 668.655 681.185 ;
        RECT 0.065 679.000 672.915 680.320 ;
        RECT 4.400 677.600 672.915 679.000 ;
        RECT 0.065 675.600 672.915 677.600 ;
        RECT 0.065 674.200 668.655 675.600 ;
        RECT 0.065 669.480 672.915 674.200 ;
        RECT 0.065 668.800 668.655 669.480 ;
        RECT 4.400 668.080 668.655 668.800 ;
        RECT 4.400 667.400 672.915 668.080 ;
        RECT 0.065 664.040 672.915 667.400 ;
        RECT 0.065 662.640 668.655 664.040 ;
        RECT 0.065 657.920 672.915 662.640 ;
        RECT 4.400 656.520 668.655 657.920 ;
        RECT 0.065 651.800 672.915 656.520 ;
        RECT 0.065 650.400 668.655 651.800 ;
        RECT 0.065 647.720 672.915 650.400 ;
        RECT 4.400 646.320 672.915 647.720 ;
        RECT 0.065 645.680 672.915 646.320 ;
        RECT 0.065 644.280 668.655 645.680 ;
        RECT 0.065 640.240 672.915 644.280 ;
        RECT 0.065 638.840 668.655 640.240 ;
        RECT 0.065 636.840 672.915 638.840 ;
        RECT 4.400 635.440 672.915 636.840 ;
        RECT 0.065 634.120 672.915 635.440 ;
        RECT 0.065 632.720 668.655 634.120 ;
        RECT 0.065 628.000 672.915 632.720 ;
        RECT 0.065 626.640 668.655 628.000 ;
        RECT 4.400 626.600 668.655 626.640 ;
        RECT 4.400 625.240 672.915 626.600 ;
        RECT 0.065 621.880 672.915 625.240 ;
        RECT 0.065 620.480 668.655 621.880 ;
        RECT 0.065 616.440 672.915 620.480 ;
        RECT 0.065 615.760 668.655 616.440 ;
        RECT 4.400 615.040 668.655 615.760 ;
        RECT 4.400 614.360 672.915 615.040 ;
        RECT 0.065 610.320 672.915 614.360 ;
        RECT 0.065 608.920 668.655 610.320 ;
        RECT 0.065 605.560 672.915 608.920 ;
        RECT 4.400 604.200 672.915 605.560 ;
        RECT 4.400 604.160 668.655 604.200 ;
        RECT 0.065 602.800 668.655 604.160 ;
        RECT 0.065 598.080 672.915 602.800 ;
        RECT 0.065 596.680 668.655 598.080 ;
        RECT 0.065 594.680 672.915 596.680 ;
        RECT 4.400 593.280 672.915 594.680 ;
        RECT 0.065 592.640 672.915 593.280 ;
        RECT 0.065 591.240 668.655 592.640 ;
        RECT 0.065 586.520 672.915 591.240 ;
        RECT 0.065 585.120 668.655 586.520 ;
        RECT 0.065 584.480 672.915 585.120 ;
        RECT 4.400 583.080 672.915 584.480 ;
        RECT 0.065 580.400 672.915 583.080 ;
        RECT 0.065 579.000 668.655 580.400 ;
        RECT 0.065 574.280 672.915 579.000 ;
        RECT 0.065 573.600 668.655 574.280 ;
        RECT 4.400 572.880 668.655 573.600 ;
        RECT 4.400 572.200 672.915 572.880 ;
        RECT 0.065 568.840 672.915 572.200 ;
        RECT 0.065 567.440 668.655 568.840 ;
        RECT 0.065 563.400 672.915 567.440 ;
        RECT 4.400 562.720 672.915 563.400 ;
        RECT 4.400 562.000 668.655 562.720 ;
        RECT 0.065 561.320 668.655 562.000 ;
        RECT 0.065 556.600 672.915 561.320 ;
        RECT 0.065 555.200 668.655 556.600 ;
        RECT 0.065 552.520 672.915 555.200 ;
        RECT 4.400 551.120 672.915 552.520 ;
        RECT 0.065 550.480 672.915 551.120 ;
        RECT 0.065 549.080 668.655 550.480 ;
        RECT 0.065 545.040 672.915 549.080 ;
        RECT 0.065 543.640 668.655 545.040 ;
        RECT 0.065 542.320 672.915 543.640 ;
        RECT 4.400 540.920 672.915 542.320 ;
        RECT 0.065 538.920 672.915 540.920 ;
        RECT 0.065 537.520 668.655 538.920 ;
        RECT 0.065 532.800 672.915 537.520 ;
        RECT 0.065 531.440 668.655 532.800 ;
        RECT 4.400 531.400 668.655 531.440 ;
        RECT 4.400 530.040 672.915 531.400 ;
        RECT 0.065 526.680 672.915 530.040 ;
        RECT 0.065 525.280 668.655 526.680 ;
        RECT 0.065 521.240 672.915 525.280 ;
        RECT 4.400 519.840 668.655 521.240 ;
        RECT 0.065 515.120 672.915 519.840 ;
        RECT 0.065 513.720 668.655 515.120 ;
        RECT 0.065 510.360 672.915 513.720 ;
        RECT 4.400 509.000 672.915 510.360 ;
        RECT 4.400 508.960 668.655 509.000 ;
        RECT 0.065 507.600 668.655 508.960 ;
        RECT 0.065 502.880 672.915 507.600 ;
        RECT 0.065 501.480 668.655 502.880 ;
        RECT 0.065 500.160 672.915 501.480 ;
        RECT 4.400 498.760 672.915 500.160 ;
        RECT 0.065 497.440 672.915 498.760 ;
        RECT 0.065 496.040 668.655 497.440 ;
        RECT 0.065 491.320 672.915 496.040 ;
        RECT 0.065 489.920 668.655 491.320 ;
        RECT 0.065 489.280 672.915 489.920 ;
        RECT 4.400 487.880 672.915 489.280 ;
        RECT 0.065 485.200 672.915 487.880 ;
        RECT 0.065 483.800 668.655 485.200 ;
        RECT 0.065 479.080 672.915 483.800 ;
        RECT 4.400 477.680 668.655 479.080 ;
        RECT 0.065 473.640 672.915 477.680 ;
        RECT 0.065 472.240 668.655 473.640 ;
        RECT 0.065 468.200 672.915 472.240 ;
        RECT 4.400 467.520 672.915 468.200 ;
        RECT 4.400 466.800 668.655 467.520 ;
        RECT 0.065 466.120 668.655 466.800 ;
        RECT 0.065 461.400 672.915 466.120 ;
        RECT 0.065 460.000 668.655 461.400 ;
        RECT 0.065 458.000 672.915 460.000 ;
        RECT 4.400 456.600 672.915 458.000 ;
        RECT 0.065 455.280 672.915 456.600 ;
        RECT 0.065 453.880 668.655 455.280 ;
        RECT 0.065 449.840 672.915 453.880 ;
        RECT 0.065 448.440 668.655 449.840 ;
        RECT 0.065 447.800 672.915 448.440 ;
        RECT 4.400 446.400 672.915 447.800 ;
        RECT 0.065 443.720 672.915 446.400 ;
        RECT 0.065 442.320 668.655 443.720 ;
        RECT 0.065 437.600 672.915 442.320 ;
        RECT 0.065 436.920 668.655 437.600 ;
        RECT 4.400 436.200 668.655 436.920 ;
        RECT 4.400 435.520 672.915 436.200 ;
        RECT 0.065 431.480 672.915 435.520 ;
        RECT 0.065 430.080 668.655 431.480 ;
        RECT 0.065 426.720 672.915 430.080 ;
        RECT 4.400 426.040 672.915 426.720 ;
        RECT 4.400 425.320 668.655 426.040 ;
        RECT 0.065 424.640 668.655 425.320 ;
        RECT 0.065 419.920 672.915 424.640 ;
        RECT 0.065 418.520 668.655 419.920 ;
        RECT 0.065 415.840 672.915 418.520 ;
        RECT 4.400 414.440 672.915 415.840 ;
        RECT 0.065 413.800 672.915 414.440 ;
        RECT 0.065 412.400 668.655 413.800 ;
        RECT 0.065 407.680 672.915 412.400 ;
        RECT 0.065 406.280 668.655 407.680 ;
        RECT 0.065 405.640 672.915 406.280 ;
        RECT 4.400 404.240 672.915 405.640 ;
        RECT 0.065 402.240 672.915 404.240 ;
        RECT 0.065 400.840 668.655 402.240 ;
        RECT 0.065 396.120 672.915 400.840 ;
        RECT 0.065 394.760 668.655 396.120 ;
        RECT 4.400 394.720 668.655 394.760 ;
        RECT 4.400 393.360 672.915 394.720 ;
        RECT 0.065 390.000 672.915 393.360 ;
        RECT 0.065 388.600 668.655 390.000 ;
        RECT 0.065 384.560 672.915 388.600 ;
        RECT 4.400 383.880 672.915 384.560 ;
        RECT 4.400 383.160 668.655 383.880 ;
        RECT 0.065 382.480 668.655 383.160 ;
        RECT 0.065 378.440 672.915 382.480 ;
        RECT 0.065 377.040 668.655 378.440 ;
        RECT 0.065 373.680 672.915 377.040 ;
        RECT 4.400 372.320 672.915 373.680 ;
        RECT 4.400 372.280 668.655 372.320 ;
        RECT 0.065 370.920 668.655 372.280 ;
        RECT 0.065 366.200 672.915 370.920 ;
        RECT 0.065 364.800 668.655 366.200 ;
        RECT 0.065 363.480 672.915 364.800 ;
        RECT 4.400 362.080 672.915 363.480 ;
        RECT 0.065 360.080 672.915 362.080 ;
        RECT 0.065 358.680 668.655 360.080 ;
        RECT 0.065 354.640 672.915 358.680 ;
        RECT 0.065 353.240 668.655 354.640 ;
        RECT 0.065 352.600 672.915 353.240 ;
        RECT 4.400 351.200 672.915 352.600 ;
        RECT 0.065 348.520 672.915 351.200 ;
        RECT 0.065 347.120 668.655 348.520 ;
        RECT 0.065 342.400 672.915 347.120 ;
        RECT 4.400 341.000 668.655 342.400 ;
        RECT 0.065 336.280 672.915 341.000 ;
        RECT 0.065 334.880 668.655 336.280 ;
        RECT 0.065 331.520 672.915 334.880 ;
        RECT 4.400 330.840 672.915 331.520 ;
        RECT 4.400 330.120 668.655 330.840 ;
        RECT 0.065 329.440 668.655 330.120 ;
        RECT 0.065 324.720 672.915 329.440 ;
        RECT 0.065 323.320 668.655 324.720 ;
        RECT 0.065 321.320 672.915 323.320 ;
        RECT 4.400 319.920 672.915 321.320 ;
        RECT 0.065 318.600 672.915 319.920 ;
        RECT 0.065 317.200 668.655 318.600 ;
        RECT 0.065 312.480 672.915 317.200 ;
        RECT 0.065 311.080 668.655 312.480 ;
        RECT 0.065 310.440 672.915 311.080 ;
        RECT 4.400 309.040 672.915 310.440 ;
        RECT 0.065 307.040 672.915 309.040 ;
        RECT 0.065 305.640 668.655 307.040 ;
        RECT 0.065 300.920 672.915 305.640 ;
        RECT 0.065 300.240 668.655 300.920 ;
        RECT 4.400 299.520 668.655 300.240 ;
        RECT 4.400 298.840 672.915 299.520 ;
        RECT 0.065 294.800 672.915 298.840 ;
        RECT 0.065 293.400 668.655 294.800 ;
        RECT 0.065 289.360 672.915 293.400 ;
        RECT 4.400 288.680 672.915 289.360 ;
        RECT 4.400 287.960 668.655 288.680 ;
        RECT 0.065 287.280 668.655 287.960 ;
        RECT 0.065 283.240 672.915 287.280 ;
        RECT 0.065 281.840 668.655 283.240 ;
        RECT 0.065 279.160 672.915 281.840 ;
        RECT 4.400 277.760 672.915 279.160 ;
        RECT 0.065 277.120 672.915 277.760 ;
        RECT 0.065 275.720 668.655 277.120 ;
        RECT 0.065 271.000 672.915 275.720 ;
        RECT 0.065 269.600 668.655 271.000 ;
        RECT 0.065 268.280 672.915 269.600 ;
        RECT 4.400 266.880 672.915 268.280 ;
        RECT 0.065 264.880 672.915 266.880 ;
        RECT 0.065 263.480 668.655 264.880 ;
        RECT 0.065 259.440 672.915 263.480 ;
        RECT 0.065 258.080 668.655 259.440 ;
        RECT 4.400 258.040 668.655 258.080 ;
        RECT 4.400 256.680 672.915 258.040 ;
        RECT 0.065 253.320 672.915 256.680 ;
        RECT 0.065 251.920 668.655 253.320 ;
        RECT 0.065 247.200 672.915 251.920 ;
        RECT 4.400 245.800 668.655 247.200 ;
        RECT 0.065 241.080 672.915 245.800 ;
        RECT 0.065 239.680 668.655 241.080 ;
        RECT 0.065 237.000 672.915 239.680 ;
        RECT 4.400 235.640 672.915 237.000 ;
        RECT 4.400 235.600 668.655 235.640 ;
        RECT 0.065 234.240 668.655 235.600 ;
        RECT 0.065 229.520 672.915 234.240 ;
        RECT 0.065 228.120 668.655 229.520 ;
        RECT 0.065 226.800 672.915 228.120 ;
        RECT 4.400 225.400 672.915 226.800 ;
        RECT 0.065 223.400 672.915 225.400 ;
        RECT 0.065 222.000 668.655 223.400 ;
        RECT 0.065 217.280 672.915 222.000 ;
        RECT 0.065 215.920 668.655 217.280 ;
        RECT 4.400 215.880 668.655 215.920 ;
        RECT 4.400 214.520 672.915 215.880 ;
        RECT 0.065 211.840 672.915 214.520 ;
        RECT 0.065 210.440 668.655 211.840 ;
        RECT 0.065 205.720 672.915 210.440 ;
        RECT 4.400 204.320 668.655 205.720 ;
        RECT 0.065 199.600 672.915 204.320 ;
        RECT 0.065 198.200 668.655 199.600 ;
        RECT 0.065 194.840 672.915 198.200 ;
        RECT 4.400 193.480 672.915 194.840 ;
        RECT 4.400 193.440 668.655 193.480 ;
        RECT 0.065 192.080 668.655 193.440 ;
        RECT 0.065 188.040 672.915 192.080 ;
        RECT 0.065 186.640 668.655 188.040 ;
        RECT 0.065 184.640 672.915 186.640 ;
        RECT 4.400 183.240 672.915 184.640 ;
        RECT 0.065 181.920 672.915 183.240 ;
        RECT 0.065 180.520 668.655 181.920 ;
        RECT 0.065 175.800 672.915 180.520 ;
        RECT 0.065 174.400 668.655 175.800 ;
        RECT 0.065 173.760 672.915 174.400 ;
        RECT 4.400 172.360 672.915 173.760 ;
        RECT 0.065 169.680 672.915 172.360 ;
        RECT 0.065 168.280 668.655 169.680 ;
        RECT 0.065 164.240 672.915 168.280 ;
        RECT 0.065 163.560 668.655 164.240 ;
        RECT 4.400 162.840 668.655 163.560 ;
        RECT 4.400 162.160 672.915 162.840 ;
        RECT 0.065 158.120 672.915 162.160 ;
        RECT 0.065 156.720 668.655 158.120 ;
        RECT 0.065 152.680 672.915 156.720 ;
        RECT 4.400 152.000 672.915 152.680 ;
        RECT 4.400 151.280 668.655 152.000 ;
        RECT 0.065 150.600 668.655 151.280 ;
        RECT 0.065 145.880 672.915 150.600 ;
        RECT 0.065 144.480 668.655 145.880 ;
        RECT 0.065 142.480 672.915 144.480 ;
        RECT 4.400 141.080 672.915 142.480 ;
        RECT 0.065 140.440 672.915 141.080 ;
        RECT 0.065 139.040 668.655 140.440 ;
        RECT 0.065 134.320 672.915 139.040 ;
        RECT 0.065 132.920 668.655 134.320 ;
        RECT 0.065 131.600 672.915 132.920 ;
        RECT 4.400 130.200 672.915 131.600 ;
        RECT 0.065 128.200 672.915 130.200 ;
        RECT 0.065 126.800 668.655 128.200 ;
        RECT 0.065 122.080 672.915 126.800 ;
        RECT 0.065 121.400 668.655 122.080 ;
        RECT 4.400 120.680 668.655 121.400 ;
        RECT 4.400 120.000 672.915 120.680 ;
        RECT 0.065 116.640 672.915 120.000 ;
        RECT 0.065 115.240 668.655 116.640 ;
        RECT 0.065 110.520 672.915 115.240 ;
        RECT 4.400 109.120 668.655 110.520 ;
        RECT 0.065 104.400 672.915 109.120 ;
        RECT 0.065 103.000 668.655 104.400 ;
        RECT 0.065 100.320 672.915 103.000 ;
        RECT 4.400 98.920 672.915 100.320 ;
        RECT 0.065 98.280 672.915 98.920 ;
        RECT 0.065 96.880 668.655 98.280 ;
        RECT 0.065 92.840 672.915 96.880 ;
        RECT 0.065 91.440 668.655 92.840 ;
        RECT 0.065 89.440 672.915 91.440 ;
        RECT 4.400 88.040 672.915 89.440 ;
        RECT 0.065 86.720 672.915 88.040 ;
        RECT 0.065 85.320 668.655 86.720 ;
        RECT 0.065 80.600 672.915 85.320 ;
        RECT 0.065 79.240 668.655 80.600 ;
        RECT 4.400 79.200 668.655 79.240 ;
        RECT 4.400 77.840 672.915 79.200 ;
        RECT 0.065 74.480 672.915 77.840 ;
        RECT 0.065 73.080 668.655 74.480 ;
        RECT 0.065 69.040 672.915 73.080 ;
        RECT 0.065 68.360 668.655 69.040 ;
        RECT 4.400 67.640 668.655 68.360 ;
        RECT 4.400 66.960 672.915 67.640 ;
        RECT 0.065 62.920 672.915 66.960 ;
        RECT 0.065 61.520 668.655 62.920 ;
        RECT 0.065 58.160 672.915 61.520 ;
        RECT 4.400 56.800 672.915 58.160 ;
        RECT 4.400 56.760 668.655 56.800 ;
        RECT 0.065 55.400 668.655 56.760 ;
        RECT 0.065 50.680 672.915 55.400 ;
        RECT 0.065 49.280 668.655 50.680 ;
        RECT 0.065 47.280 672.915 49.280 ;
        RECT 4.400 45.880 672.915 47.280 ;
        RECT 0.065 45.240 672.915 45.880 ;
        RECT 0.065 43.840 668.655 45.240 ;
        RECT 0.065 39.120 672.915 43.840 ;
        RECT 0.065 37.720 668.655 39.120 ;
        RECT 0.065 37.080 672.915 37.720 ;
        RECT 4.400 35.680 672.915 37.080 ;
        RECT 0.065 33.000 672.915 35.680 ;
        RECT 0.065 31.600 668.655 33.000 ;
        RECT 0.065 26.880 672.915 31.600 ;
        RECT 0.065 26.200 668.655 26.880 ;
        RECT 4.400 25.480 668.655 26.200 ;
        RECT 4.400 24.800 672.915 25.480 ;
        RECT 0.065 21.440 672.915 24.800 ;
        RECT 0.065 20.040 668.655 21.440 ;
        RECT 0.065 16.000 672.915 20.040 ;
        RECT 4.400 15.320 672.915 16.000 ;
        RECT 4.400 14.600 668.655 15.320 ;
        RECT 0.065 13.920 668.655 14.600 ;
        RECT 0.065 9.200 672.915 13.920 ;
        RECT 0.065 7.800 668.655 9.200 ;
        RECT 0.065 5.800 672.915 7.800 ;
        RECT 4.400 4.400 672.915 5.800 ;
        RECT 0.065 3.760 672.915 4.400 ;
        RECT 0.065 2.360 668.655 3.760 ;
        RECT 0.065 0.175 672.915 2.360 ;
      LAYER met4 ;
        RECT 0.295 672.480 663.025 679.825 ;
        RECT 0.295 10.240 20.640 672.480 ;
        RECT 23.040 672.240 97.440 672.480 ;
        RECT 23.040 10.480 23.940 672.240 ;
        RECT 26.340 10.480 27.240 672.240 ;
        RECT 29.640 10.480 30.540 672.240 ;
        RECT 32.940 10.480 97.440 672.240 ;
        RECT 23.040 10.240 97.440 10.480 ;
        RECT 99.840 672.240 174.240 672.480 ;
        RECT 99.840 10.480 100.740 672.240 ;
        RECT 103.140 10.480 104.040 672.240 ;
        RECT 106.440 10.480 107.340 672.240 ;
        RECT 109.740 10.480 174.240 672.240 ;
        RECT 99.840 10.240 174.240 10.480 ;
        RECT 176.640 672.240 251.040 672.480 ;
        RECT 176.640 10.480 177.540 672.240 ;
        RECT 179.940 10.480 180.840 672.240 ;
        RECT 183.240 10.480 184.140 672.240 ;
        RECT 186.540 10.480 251.040 672.240 ;
        RECT 176.640 10.240 251.040 10.480 ;
        RECT 253.440 672.240 327.840 672.480 ;
        RECT 253.440 10.480 254.340 672.240 ;
        RECT 256.740 10.480 257.640 672.240 ;
        RECT 260.040 10.480 260.940 672.240 ;
        RECT 263.340 10.480 327.840 672.240 ;
        RECT 253.440 10.240 327.840 10.480 ;
        RECT 330.240 672.240 404.640 672.480 ;
        RECT 330.240 10.480 331.140 672.240 ;
        RECT 333.540 10.480 334.440 672.240 ;
        RECT 336.840 10.480 337.740 672.240 ;
        RECT 340.140 10.480 404.640 672.240 ;
        RECT 330.240 10.240 404.640 10.480 ;
        RECT 407.040 672.240 481.440 672.480 ;
        RECT 407.040 10.480 407.940 672.240 ;
        RECT 410.340 10.480 411.240 672.240 ;
        RECT 413.640 10.480 414.540 672.240 ;
        RECT 416.940 10.480 481.440 672.240 ;
        RECT 407.040 10.240 481.440 10.480 ;
        RECT 483.840 672.240 558.240 672.480 ;
        RECT 483.840 10.480 484.740 672.240 ;
        RECT 487.140 10.480 488.040 672.240 ;
        RECT 490.440 10.480 491.340 672.240 ;
        RECT 493.740 10.480 558.240 672.240 ;
        RECT 483.840 10.240 558.240 10.480 ;
        RECT 560.640 672.240 635.040 672.480 ;
        RECT 560.640 10.480 561.540 672.240 ;
        RECT 563.940 10.480 564.840 672.240 ;
        RECT 567.240 10.480 568.140 672.240 ;
        RECT 570.540 10.480 635.040 672.240 ;
        RECT 560.640 10.240 635.040 10.480 ;
        RECT 637.440 672.240 663.025 672.480 ;
        RECT 637.440 10.480 638.340 672.240 ;
        RECT 640.740 10.480 641.640 672.240 ;
        RECT 644.040 10.480 644.940 672.240 ;
        RECT 647.340 10.480 663.025 672.240 ;
        RECT 637.440 10.240 663.025 10.480 ;
        RECT 0.295 0.175 663.025 10.240 ;
      LAYER met5 ;
        RECT 33.700 269.600 382.140 305.100 ;
        RECT 33.700 193.010 382.140 254.660 ;
        RECT 33.700 116.420 382.140 178.070 ;
        RECT 33.700 39.830 382.140 101.480 ;
        RECT 33.700 0.900 382.140 24.890 ;
  END
END wrapper_sha1
END LIBRARY

