module dump();
    initial begin
        $dumpfile ("wrapper.vcd");
        $dumpvars (0, wrapper_sha1);
        #1;
    end
endmodule
